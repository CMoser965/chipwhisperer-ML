module parameters (
	output logic [31:0][0:0][8:0] weights_o_0,
	output logic [31:0][2:0] threshold_o_0,
	output logic [31:0][1:0] sign_o_0,
	output logic [287:0][63:0] weights_o_1,
	output logic [63:0][9:0] threshold_o_1,
	output logic [63:0][1:0] sign_o_1,
	output logic [0:0][63:0][9:0] weights_o_2,
	output logic [9:0][4:0] threshold_o_2,
	output logic [9:0][1:0] sign_o_2
);

// assign weights
assign weight_o_0 = {{9'b010010010},{9'b001111001},{9'b011001000},{9'b001101011},{9'b100110001},{9'b010000100},{9'b000100001},{9'b000111101},{9'b000010011},{9'b100110001},{9'b000000111},{9'b000100001},{9'b010000101},{9'b000000110},{9'b110011010},{9'b010111100},{9'b111011001},{9'b110101100},{9'b100000001},{9'b110101010},{9'b110011111},{9'b100100100},{9'b100111000},{9'b101010110},{9'b001100000},{9'b000001011},{9'b110101101},{9'b000110000},{9'b011101000},{9'b011010111},{9'b000001001},{9'b101010110}};
assign weight_o_1 = {{64'b0011110101001010011111111001111011010100101101100011011110111000},{64'b0010110000000110100010110001010111001100011111011000000010110010},{64'b1100001010110001010101001110100100000011010000101101101101111101},{64'b0011111101010010001011111001101101110000101110001101010010110000},{64'b0011010110011110110110110000001111010111101011011111011011011111},{64'b1000111111100001011101011111110000111010010010111001101100000111},{64'b1101001011010001000000010111001010000011010000100000001001110011},{64'b1100111000001001111110110010110001000000011011011111001101101100},{64'b0011010101011110011010111001110111111100001010001110010010110000},{64'b0011000001001010010010111001011011010101101101001100000010110001},{64'b0000111110110010000111010110010000100000010010111001111111100011},{64'b0101110000100011100100010111000010000000010110011100101110110010},{64'b1111001101011001111011101101010101111010101001000001100110001011},{64'b0111000001010011010101000011110111000011001100101100011111111001},{64'b1100001011110001011101001110100100100010010000101101101101001001},{64'b0101010110011110011111001111001100010101110110111100011100110110},{64'b0011110110110110101110110100001011111100000011010110000011000110},{64'b0010111100100110100100110011101100111100011111011111011000101100},{64'b1000111010101111001010010100011000101100110110101011101111000000},{64'b0010010010000010010001110001110000000100110100011100000110000000},{64'b1100001011110001001001011110101000000011110000110011101100001100},{64'b1000101110100111101100001110101000101010110110111111111000011110},{64'b1100001011110001001100110110001010100111010100011000101001011011},{64'b0011110001001010000000110001011011000101011110001000000110110011},{64'b1100101010100001011001001110110000100010110000110011101100001100},{64'b1011011001110001011001111011110101110000001110000000000010110001},{64'b1100011111110001011101011110110000000011010101111000101111001101},{64'b0011110100011100101010110000011111111101001110001100000010100011},{64'b1100001010110001001101001110100000100011110000100011101101001100},{64'b0010110000101110000011110001011011001100011111011100000110110000},{64'b1111000001000000010000101000110111110111101100000001110011111011},{64'b0111010101001010010011110011010111000001001100001100010111110011},{64'b0011001101010010011001101001101111110001101100001101000010110011},{64'b0011001001010110001111001011101111110001101110101111000010110110},{64'b0110001010110001101100100110001110001001010000011111101000001111},{64'b0010001100110110011001101001101101111011101110001111010011110100},{64'b0011100010011111001100100010101111010101111100000111110011011111},{64'b0011111011110111101000111111101101111011101000001111001010010111},{64'b0100110011111001000000110110111010100111010100011000100010000011},{64'b0010110010011110100101000010100110101110011010101111110000001001},{64'b0011010001011110111111000011100111110001101010001111001011110011},{64'b1011001001100110111010101101001001111011101011010110001000110111},{64'b1011100100101101111110101100001010011101100001010001110011001111},{64'b1100111010111010010010010110011000001110010001111000101100001111},{64'b1101001011101101110111000110110100000011010000110111101101001011},{64'b1100001010100111110101001110001000110011110010111111101101011101},{64'b1010110010100001100101010110100110000010010010101111101000001001},{64'b0011010011000110000110001000001111110111111110111110011011110111},{64'b0010101100110110001000101001101101111101101011001111011000110110},{64'b0100101100110010011001111111101000011010100101011111011100110100},{64'b1000101010111111111010100100001000111111101011000111100000011111},{64'b0011101000011110101100101000001111011101101010000111010000100100},{64'b1100001010110001000000010110010010001110010101110001101101001111},{64'b0010100010111101001000100000001011101101011111010000100010000111},{64'b0101000010001110000100010010111010000101010101101000001001011000},{64'b0011000111010110010110101000001111010101101110001111010011110101},{64'b1100101001110001001001110110011010101011010100000001100011011110},{64'b1100101010100111111110001110001000101011110010111111101100001101},{64'b0000110010001000010010110100011010101100010111011000100110001111},{64'b0111001001011111110110000011101111000011101000101100011111110011},{64'b1100101010110001001000110110010010001011010100000001101000001111},{64'b0011010110011110110100001100101001111101100111101111110111111100},{64'b1000111010110111111110001100011000111110110011110011111100001100},{64'b1101000011011101110111000110100100000011000010110110000001110001},{64'b1100111011101110110111011111101000110010100010111110001101110001},{64'b1110011101100010111111011111100101110010101000100111011100110000},{64'b0011000000010011001000100000000111011101001101000001010011111110},{64'b1101011101101110010001011111101100010011100110101111011111110100},{64'b0000101110110010001000101100001110111111101111001111110010110111},{64'b0001000001001111001100001010010111010110110100100011011011111100},{64'b1100111010100100010101011110011000101010010011111010101100000101},{64'b0000101110110010001000101000001111111110100101001001010011110110},{64'b1111010101001111110111011011100101000011101010101100001101110001},{64'b1101011000100101111111011111101000110011100011111110011100010001},{64'b0101000101001010011001111001110111000100000101000000000111110010},{64'b1011001001011000101000100100010010000101010001100000101011000111},{64'b1011000010101101110110010110001000100001111011111110101100010001},{64'b1000111010101101101010010110001000101011110011111010101100000111},{64'b0010110010110010001000100001111110110110101100101001010011110110},{64'b1101011001101101110111011111100000000010110011111110111100010001},{64'b1111010101001110110111001011110101000011001010100100001101111000},{64'b1100111111110010111011001111110001111010100010110001100110000001},{64'b0001000001001101100110110010010010001101010001000000101111001011},{64'b0010110100110010000000111001111111110100001101001001010011110110},{64'b1110001100010001001000100000001111111110101101000001110010101110},{64'b0101000101011111011110001100011111010111101101100001110011111110},{64'b0100101010110011000000111110011010011111110101011011110000010100},{64'b0110001101010010001001111001110111010101101100001101000011110110},{64'b0010000010010000001000101100001110011110111101000001110011111110},{64'b1011000000101101110110110110001010001001101011111110101100000011},{64'b0001010000001001110111110000010001000100010110000000100111100100},{64'b1101001010101101110111011110101000000011110010111110101101010001},{64'b0110001001010001001000100000010111111100011101000001100011001110},{64'b0111000101001011011111000011110111010011001100100101000111111000},{64'b1001101010100101100000110110001010001011110011111110001000010011},{64'b0001010001001001100000110000010010000101010101001000101110000011},{64'b0100001011110010011000111011001011110011101010001100001000110111},{64'b1011111010110100101100010110000100011000011110101101111000100010},{64'b0000110101001110110110000001010111000100010100110000110111001000},{64'b0111001001100110010000110011001011010001101110001110000110110111},{64'b1100101011111001011001001100010110100111000000100001100111001111},{64'b0101011101101100110011111001111000000100000001111000001101010000},{64'b0001010010001101100111000010110101100000000010111111110001001000},{64'b1100001011110001010001011110110110100011010100101001100011001011},{64'b0111000100101110000010101010011010010101100111011110011111010110},{64'b1001011001100011110101011011100101000010001000101111111001101010},{64'b1111001001110001011101011111100000100011011000101111101000011011},{64'b0111111010000111001101010011000111000011011110101111011001011111},{64'b0011110101001110111010111001011101111100001111010010010111110100},{64'b0001110101001110110010010101010001011000100111010010010111100100},{64'b0000110101001010110011000101110110000100010101100000110111101000},{64'b1100101111000001101100111100000000101011010010010011101100001011},{64'b0011010100001100111011110001010011011100101011011110001100110000},{64'b0111001011010011000000110011001010010011101100001100000010110111},{64'b1101001001111001001001110011000010000011001000101110001000010011},{64'b1110101011110001011001011111110010100011011000101000100100010011},{64'b0000000110001101110101001010010111000110010100101011110101101000},{64'b0001000011001101110000100000010111000110000100000100010001001001},{64'b1110110011010001110101000110110110100010011000100001110001001011},{64'b0100001001110001001101010011110111100010011100100101001100001010},{64'b1100000100001010110000001011110110001110000101111011110101101000},{64'b0001100100001100000010100001111001000100001101011010011111110000},{64'b1101001001111001010101001111100100000011000000101111111000001001},{64'b0011111010010110100100100000101111010001011110101111011001011111},{64'b1001010110001110010010000100111111000100000100110011110111101000},{64'b0001101110000100101101010001100100111000011011110111001000101000},{64'b0011110101101110110110011101001101111000101111010010010111110000},{64'b0001011110101100110111000101110000000000100111111010111101011010},{64'b0011001011010101101000101000001111011001101001000101010010010111},{64'b0110001001000010001000110010001110010101100100001000001011110110},{64'b0101000100001101110010001000011110000110100101110011110001001100},{64'b0011001011101111001100000110001000110001101000101100001000110011},{64'b0110000010010001000000100010001110000111010100101001000011011111},{64'b1100001100101101001100001110111010011011100001110011111101011100},{64'b1011010101000000100101110011100101100000001010001110001000111000},{64'b0011000010111010000000110010011110010101111100001001010011110110},{64'b0011001010110010001000001000001011111101101101100101001011011110},{64'b0011010000000100100101110011100100000000001110001110011100111000},{64'b1110111101110010000101111101101001111010011110101100100110100011},{64'b0000110110000000110111001101110101100110000101111011110111101000},{64'b1101000101101101110010000101010000001000100011110000010101000001},{64'b1011110100001100111111100001110111111100001111010011110011101000},{64'b0101001001001110010000010010101010000011110100101000010101010111},{64'b0111011001110001101101010010100110010011101100101100011000111011},{64'b1101001011110011010100010110001000110011110000101100101010010111},{64'b0100110011101100111010110011001010001001010011010000100110000001},{64'b1010110110010110110111011101110101110100011110001010110110100000},{64'b0110001011110011000000110010001010010111011100101101100011011111},{64'b1100000100001001110010001001110101000110010101110011110111001000},{64'b1100011011100001111111001111110000000011110000110000101100001000},{64'b1010111010100101100101010110100101100010011010101110100010001011},{64'b0111001011010001001100100110001000010011001010101111101010010111},{64'b1100000100001001111001001010110001001110100101110011111101001100},{64'b1100000101001011010011101111110000000110100101110000110111001100},{64'b1010111101110000101011111101100101110000011110001010100110100001},{64'b0011010000110110000101010011100110110001101110001110011010110011},{64'b1101000100001101110010001110110100000100000001111010110111001000},{64'b1111001011110110010100011110001001110011111110101110100010010011},{64'b1100010101101000110001101001110101000000100001010011010101100000},{64'b0100000100001101101101101010110100000100011001110111110001001000},{64'b1001110011011111110111010101010101100010010110100000100111001001},{64'b1101110011100110110111010110101000000010010010111110101101011001},{64'b1101111111001111110111010111010001100011010010111100101110000001},{64'b0101111011101110110110010111001010000001100010111100001100110001},{64'b1000111111111001111110101100010011111001010001010001100111000111},{64'b1011001111011111111110001110001111111011101010110111011001010011},{64'b0010010010010110000001011010110111000100011100100111110011101100},{64'b1010100100011001011110101101010111101100011101000001110011001110},{64'b0011000011001111100100110010001010001101101010011110001001110011},{64'b1011000000010001101101101001100111110010001100000101110001101110},{64'b0010111010100110000000010000101100010001011011111110011110001010},{64'b0000010100110010010000101101101100110110101101101011110010111100},{64'b0101001001101101111000111011001010010001101011010110001000010111},{64'b0000001000110110011000100101001100011101100111000011010111110100},{64'b0011000101011001001000100001010111111101101001010000110111001010},{64'b1011000000010101100111000000100101110010101000100111111011101000},{64'b0001011001101110110010010110001000000001100011111110001100110001},{64'b0100100100110000001001101100011010111101011101011000100110001110},{64'b1110101100010001011001111101111111110100101101010001110110101110},{64'b1110100100011001011001100001010111101100011001000001110111001010},{64'b0010110001011011010010111111101001100101001110001110110010100011},{64'b1101111111100011110111011101011001101000000010011000000110110011},{64'b1110101010010001001001001010100111010110111100100001110001101110},{64'b1100111110100000110001111110110000101000010001111000100100001000},{64'b1011001011010111001100001001001101110111101010000111110011011011},{64'b0011000000101110101010101000001101111001101011011110000000010111},{64'b0010000100000100000001110001110101010100101101001011010011100000},{64'b0010100110010010001000101000001110011101111101000111110011001110},{64'b0001111111011111010110010101001000100000000010101000110110110011},{64'b1001011001101110111010011110001000110001101011111110001000010101},{64'b1100000101101101011001101110001001011111100010010111111100010101},{64'b1110101100010001001001101001110101111000101101000001010110101010},{64'b1110011011010011010101010111100110100011011010101100101000110011},{64'b0000011111111011010110011100011001110001010110101000100110010111},{64'b1010100100000001101011110001100001001000101011010011111000001010},{64'b1011101011100011000110110010000000110011011010001100000000110011},{64'b0101100010010110000100010110111100010110010100011111011101111110},{64'b1000110010011011010110111101000001111000011111010000101000101001},{64'b0001000100001100101001001000110101000000101001010111011101111100},{64'b0000110110100110000100000000111100001100010101101011011101111100},{64'b1011111111111010011111010110001010111000011011100010000110010011},{64'b1100011111001111110011001110011101001010000010101101111111010100},{64'b1100001110111111100100001110110110001111000100100001111001001100},{64'b1100000100001101111010000100110110001110100001010001110001001100},{64'b1010111001110001001011110101100001111000101011001100000010110011},{64'b0101000100001100111000101010111000001000101001010110011101111100},{64'b0011110101000100100111110001000001101000011011011110001110100010},{64'b0100011010110010010001011100111000010011100100101110010111110100},{64'b1011111011110010010011111111001001110001101110001100000110110011},{64'b0011001010011111100100000000001111111011011110101101010011011001},{64'b1100001010000011111000001010100110001111110000110001110001001100},{64'b0100010010001110000101010010110110000000010100111111111101101100},{64'b1110110100001101111010001100010101101100000111010001111111001010},{64'b1011111001110001101111111011100111110000111010000101001000101011},{64'b0100000100000010110001001000110101010000100101110011111101101100},{64'b1100010100111011011001001100110100011110100100100001111101001100},{64'b0110110100001101110010100001110111001100001101100011100101001000},{64'b0010010000110011101001110001001111111000011101000010101010001110},{64'b1100000100001001101101001100110111001110000001100001111001001100},{64'b1010111011110011010110000100001111111011010110101101100110000011},{64'b1000100100000101101011100101100110101000000011010010101100001000},{64'b1010111111111011111110100101011001111110001010100001100010001001},{64'b0111001000101101101000101010001010010001101011011110001000110111},{64'b1101000100001001111001101000110101000010100001010011111101001100},{64'b1010111010110000001101110111001110101111011010001100000010001011},{64'b0101000011011110010110000100011011010111010100101100000111110101},{64'b1011110010110110101111111010101101111000101011000111000010110011},{64'b0101000111011110010110001100011101100111000100100100110111110101},{64'b0001000011010110000110001010101101110011110100101111011011110101},{64'b0101000000001111110100010010011010000111100100111110010101010100},{64'b1011001000000101101101100011000111101001101011001101011000101011},{64'b0011010010000110100100010010101100010000111110101111011001110100},{64'b0100010011111110010110010100011100010111010110101000100111110101},{64'b0001000000000001101101000010100110001110100001100111011001001100},{64'b0101000000001001001000101010100010000111100001010001111001011110},{64'b1110001100111001101001101011101011011011101001010101101000001111},{64'b0011011000100110001111010001101110010111001110111110011101110010},{64'b1011001001111101101100101011001001111011101010010111001010010111},{64'b0011110010100110100100010011101110111011011010111111001001101100},{64'b0101000010001111100000000010011110000011110110111110011001010101},{64'b0101000011001110010110010110111100000111010100101110010111110100},{64'b0011100001110110000000101011111000110000111011001011000011111110},{64'b0110001100110001001000101010001110011111101101010001101001001110},{64'b0011110110000110100110001000110100000110000111101111111111001100},{64'b1010101100000001101001101011110011101000001001010001101000001110},{64'b1101001000101101001000101010100110111111100001010011111000011111},{64'b0011010100000100101101000000100101001100101110101111011001111100},{64'b0101000011011101001100100010001110010111101000000011100001011111},{64'b1111010100001101111011111001100001101000101011010100001100001010},{64'b1011011101110110001011001001101101110010001110100111010011110110},{64'b0111001000001001001000101010110010001111101001010101011001011110},{64'b0011000000011101000000100010101110000111101100101110010011110110},{64'b1010110100000001101001101011110011101100001011010001101000101010},{64'b0000001011111011010000000110011010010111110100100001100011001101},{64'b1011111101110001001101111011101001111001111011000101001000110011},{64'b0011000010011111101100000000001111011111111110101101101011011111},{64'b0100111001101010011001111011111000000000100101011100001100110000},{64'b0100000101001110010010101001011011001101100101010000010111110100},{64'b1010101000100001001001111011101010111001101011011111001000101111},{64'b0101000100001101101000101000010011001101101001010000001101000110},{64'b0111000000011110010001111010111101010011101100101111011011110111},{64'b0101000111001110010100100100011111110111101100110110010011110111},{64'b1110101111011101101110001101000001101010000010100001111101001011},{64'b0001000000010010000101110010111100000011101100101111010000111101},{64'b0101000111011110110110000100011001000101010101110000110111010110},{64'b0101111101010100101010010001101001001010010010111000011110110001},{64'b1110110100001001101011100100110011101000001011010001101000001010},{64'b1010111110000001111111010011000101111010011010101111000000101000},{64'b1010110010110100100101010110100101111010011010101101101000001011},{64'b1100010110011110110110001100110111000110010001110011111001011100},{64'b1110001010110000000101010010100100100010110000111111011000111000},{64'b0011000001101101110110110000011011011101011111000100000011010011},{64'b1011110010000000100100100000100111111101011111010101111010001001},{64'b1110010101100001111111101101100001110010001010000110110000000001},{64'b1010111010110011101100000100100110110010010010101101101000101011},{64'b0100001000010010000001110010101110000011101100001111000100110110},{64'b1110111101100001011111001101100101110010011000000101100010101000},{64'b0111001100101100001000101000101010011001101001010111010000110110},{64'b1010111010010001101101010010100100111010011010101101111000001011},{64'b0101001100000010001000111010111010011101100101001001001111110100},{64'b1001111110111111010110100111001000010110011101100001000011111111},{64'b0001010111001100111110010000011011001101010011010000101011000010},{64'b0010001010100101101101101010100110010110101000011101011000101111},{64'b1101101101011001111011101101010101111010101001110001110111000011},{64'b1010111100000001101100101011101111111000101011011110011010101100},{64'b0111000000001101101000100000111111001101001101000001010011011110},{64'b0101010110100110100110001000010110011000110111100111111011111100},{64'b1010110010110110100101010110100110101110010110101101101000001001}};
assign weight_o_2 = {{10'b0111000110},{10'b1001101100},{10'b1110110010},{10'b1101110000},{10'b0010001011},{10'b1010101011},{10'b1101001110},{10'b0101001011},{10'b0110010101},{10'b0100100110},{10'b0011001111},{10'b0110011110},{10'b1101110010},{10'b1100100001},{10'b0100101101},{10'b1110010110},{10'b1100110011},{10'b0101100110},{10'b0101011010},{10'b0110110000},{10'b1100100011},{10'b0011101110},{10'b1000011010},{10'b1010001111},{10'b1101001011},{10'b0111000011},{10'b1011100110},{10'b0000101110},{10'b0011101100},{10'b0001010110},{10'b1100001101},{10'b0111111000},{10'b1100010100},{10'b0100111010},{10'b0110001010},{10'b0100001101},{10'b1101001001},{10'b0010010001},{10'b0111101100},{10'b1100000110},{10'b1101001000},{10'b0010011111},{10'b1110110010},{10'b0010111101},{10'b1110101011},{10'b1001011011},{10'b0111100001},{10'b1001001011},{10'b1010101100},{10'b1110100000},{10'b1101000001},{10'b0111011000},{10'b0110010111},{10'b0101011001},{10'b1011100001},{10'b0001100110},{10'b0100011111},{10'b0101110001},{10'b0011101000},{10'b1100101101},{10'b0011110000},{10'b1001001101},{10'b0010010110},{10'b1110000110}};
// assign threshold
assign threshold_o_0 = {3'd1,3'd2,3'd1,3'd3,3'd3,3'd3,3'd1,3'd3,3'd4,3'd1,3'd1,3'd0,3'd0,3'd1,3'd2,3'd2,3'd2,3'd1,3'd1,3'd2,3'd2,3'd1,3'd4,3'd2,3'd3,3'd1,3'd1,3'd3,3'd1,3'd3,3'd0,3'd2};
assign threshold_o_1 = {10'd228,10'd562,10'd614,10'd456,10'd201,10'd65,10'd401,10'd375,10'd232,10'd294,10'd544,10'd29,10'd719,10'd230,10'd64,10'd710,10'd380,10'd168,10'd435,10'd415,10'd326,10'd54,10'd247,10'd440,10'd308,10'd239,10'd77,10'd590,10'd188,10'd328,10'd26,10'd38,10'd467,10'd107,10'd275,10'd705,10'd498,10'd674,10'd189,10'd433,10'd146,10'd372,10'd636,10'd23,10'd308,10'd144,10'd308,10'd254,10'd274,10'd76,10'd469,10'd99,10'd557,10'd286,10'd347,10'd44,10'd313,10'd221,10'd942,10'd17,10'd331,10'd383,10'd491,10'd22};
assign threshold_o_2 = {5'd13,5'd16,5'd3,5'd7,5'd1,5'd19,5'd10,5'd10,5'd10,5'd3};

// assign sign
assign sign_o_0 = {2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd0, 2'd0, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd0, 2'd1};
assign sign_o_1 = {2'd1, 2'd1, 2'd0, 2'd1, 2'd1, 2'd1, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd0, 2'd0, 2'd0, 2'd1, 2'd1, 2'd1, 2'd1, 2'd0, 2'd1, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd1, 2'd0, 2'd1, 2'd1, 2'd1, 2'd1, 2'd0, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd0, 2'd1, 2'd0, 2'd0, 2'd0, 2'd1, 2'd0, 2'd0, 2'd0, 2'd0, 2'd0, 2'd0, 2'd1, 2'd0, 2'd0, 2'd0, 2'd1, 2'd0, 2'd1, 2'd0, 2'd0, 2'd0};
assign sign_o_2 = {2'd1, 2'd0, 2'd1, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd1, 2'd1};
endmodule

