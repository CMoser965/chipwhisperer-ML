module stimulus();

logic [27:0][27:0] mem_image;
logic [2:0][2:0] kernel;
logic clk = 1'b1;

initial begin
    mem_image[0] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[1] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[2] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[3] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[4] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[5] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[6] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[7] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[8] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[9] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[10] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[11] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[12] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[13] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[14] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[15] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[16] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[17] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[18] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[19] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[20] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[21] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[22] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[23] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[24] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[25] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[26] = 28'b1010_1010_1010_1010_1010_1010_1010;
    mem_image[27] = 28'b1010_1010_1010_1010_1010_1010_1010;
    kernel[0] = 3'b101;
    kernel[1] = 3'b010;
    kernel[2] = 3'b101;
end

logic [25:0][25:0][3:0] output_image;

BConv_Interface DUT(
    .layer_i(mem_image),
    .kernel(kernel),
    .clk(clk),
    .layer_o(output_image)
);

always #5 clk = ~clk;

initial begin
    // #1000 clk =1'b0;
    // #2000 $finish();
end

endmodule