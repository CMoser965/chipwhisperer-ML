module stimulus();



endmodule