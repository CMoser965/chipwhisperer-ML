module parameters (
	output logic [31:0][0:0][8:0] weights_o_0,
	output logic [31:0][3:0] threshold_o_0,
	output logic [31:0][1:0] sign_o_0,
	output logic [63:0][31:0][8:0] weights_o_1,
	output logic [62:0][8:0] threshold_o_1,
	output logic [63:0][1:0] sign_o_1,
	output logic [575:0][63:0][8:0] weights_o_2,
	output logic [575:0][9:0] threshold_o_2,
	output logic [575:0][1:0] sign_o_2,
	output logic [63:0][575:0] weights_o_4,
	output logic [63:0][10:0] threshold_o_4,
	output logic [63:0][1:0] sign_o_4,
	output logic [9:0][63:0] weights_o_5
);

// assign weights
assign weight_o_0 = {{9'b100111101}, {9'b110000010}, {9'b110100100}, {9'b010000010}, {9'b100010001}, {9'b000111001}, {9'b000001100}, {9'b101101010}, {9'b000000001}, {9'b110100000}, {9'b010101010}, {9'b011100101}, {9'b011101000}, {9'b010111010}, {9'b000100000}, {9'b001000101}, {9'b111000001}, {9'b100100001}, {9'b110010000}, {9'b101000110}, {9'b000101110}, {9'b011010011}, {9'b111101011}, {9'b110001011}, {9'b111110100}, {9'b100100111}, {9'b010111110}, {9'b011011100}, {9'b011011110}, {9'b011101101}, {9'b011101010}, {9'b101000011}};
assign weight_o_1 = {{9'b000010000},{9'b100000000},{9'b010000101},{9'b111010011},{9'b101000000},{9'b010111001},{9'b001000111},{9'b110101001},{9'b100011000},{9'b100011011},{9'b010100001},{9'b001110001},{9'b100111000},{9'b000110011},{9'b000110111},{9'b101000000},{9'b110000001},{9'b001101010},{9'b011101111},{9'b000001100},{9'b011001100},{9'b110000011},{9'b001111010},{9'b001001010},{9'b100101000},{9'b010111101},{9'b010010111},{9'b101100000},{9'b111110001},{9'b011101101},{9'b011111010},{9'b111111101},{9'b111101011},{9'b001101100},{9'b000101110},{9'b110001001},{9'b101110000},{9'b100011111},{9'b100001010},{9'b011100111},{9'b000010101},{9'b011001001},{9'b001011000},{9'b010111111},{9'b110000100},{9'b111101100},{9'b000010011},{9'b100011011},{9'b000111101},{9'b101000101},{9'b011100111},{9'b110001000},{9'b000101001},{9'b011010110},{9'b011100111},{9'b010110101},{9'b111001010},{9'b000101010},{9'b010100101},{9'b100111110},{9'b110011110},{9'b001100110},{9'b010010010},{9'b110001101},{9'b100010111},{9'b011010010},{9'b110111010},{9'b001011111},{9'b000010010},{9'b111001001},{9'b011100110},{9'b110010100},{9'b010100001},{9'b000000000},{9'b001011100},{9'b110100100},{9'b011001101},{9'b111000001},{9'b010011100},{9'b111100101},{9'b101010100},{9'b001000111},{9'b011000100},{9'b101101010},{9'b101010000},{9'b101111110},{9'b100100001},{9'b011000001},{9'b000010111},{9'b001011011},{9'b100100001},{9'b010010010},{9'b001001011},{9'b000111011},{9'b000101100},{9'b011010100},{9'b100011110},{9'b101001111},{9'b110000110},{9'b011000000},{9'b101111111},{9'b111011101},{9'b010100010},{9'b011011000},{9'b000100110},{9'b010110111},{9'b100101101},{9'b010001110},{9'b011011010},{9'b011100101},{9'b011111100},{9'b000011010},{9'b100000111},{9'b000110010},{9'b101001001},{9'b010010010},{9'b000011111},{9'b100011001},{9'b000001000},{9'b110001000},{9'b110001001},{9'b110100101},{9'b101111101},{9'b000101111},{9'b000000101},{9'b111100010},{9'b110100100},{9'b010010000},{9'b111010110},{9'b010111000},{9'b110011101},{9'b110110010},{9'b010110111},{9'b001000001},{9'b000101100},{9'b010010100},{9'b111100101},{9'b000010101},{9'b000011000},{9'b100100100},{9'b011011101},{9'b110100001},{9'b101101111},{9'b111000101},{9'b111110010},{9'b101101110},{9'b011001101},{9'b001001010},{9'b111010101},{9'b111001110},{9'b001100000},{9'b010000000},{9'b011100010},{9'b001101101},{9'b000111010},{9'b011001100},{9'b111001000},{9'b110110101},{9'b110100101},{9'b101000110},{9'b110110101},{9'b110111010},{9'b110111011},{9'b011110100},{9'b100011111},{9'b101111010},{9'b100101000},{9'b010011011},{9'b010101101},{9'b111111010},{9'b001111110},{9'b011111010},{9'b110001010},{9'b110111001},{9'b001111001},{9'b000000111},{9'b001001010},{9'b100110101},{9'b101010101},{9'b111100110},{9'b101011010},{9'b000011000},{9'b110001101},{9'b010110000},{9'b100111111},{9'b010110010},{9'b101110111},{9'b111110100},{9'b111011100},{9'b000000110},{9'b101011001},{9'b111101100},{9'b110011110},{9'b101010011},{9'b010111001},{9'b011101011},{9'b000110110},{9'b101000011},{9'b000010101},{9'b010101010},{9'b100011000},{9'b111111010},{9'b100100011},{9'b101101001},{9'b101100100},{9'b010010011},{9'b010101110},{9'b001110101},{9'b001101010},{9'b001101010},{9'b011011011},{9'b101101010},{9'b001010111},{9'b111100011},{9'b001111110},{9'b000101000},{9'b010101110},{9'b001101111},{9'b010110111},{9'b101101010},{9'b110100101},{9'b111110000},{9'b001110101},{9'b011111010},{9'b001011010},{9'b011100111},{9'b110011011},{9'b100100001},{9'b011101010},{9'b000100000},{9'b101010100},{9'b110110111},{9'b010111110},{9'b110101100},{9'b101110111},{9'b010010011},{9'b100000111},{9'b010111101},{9'b000010111},{9'b100011011},{9'b110011001},{9'b001111011},{9'b101111000},{9'b001011000},{9'b011010100},{9'b010101101},{9'b001011100},{9'b011000111},{9'b011010001},{9'b100101100},{9'b011100110},{9'b110111101},{9'b110000010},{9'b110010101},{9'b101110111},{9'b101001010},{9'b011011110},{9'b110101111},{9'b100101111},{9'b011110011},{9'b110110011},{9'b011001110},{9'b001001000},{9'b101010010},{9'b111000110},{9'b000101011},{9'b010100010},{9'b110000100},{9'b001000111},{9'b001010101},{9'b011100110},{9'b101101110},{9'b010010101},{9'b011010001},{9'b001101011},{9'b110001100},{9'b110101001},{9'b010001111},{9'b001100000},{9'b110111010},{9'b000011011},{9'b101000010},{9'b001000101},{9'b101110001},{9'b010100101},{9'b011010101},{9'b010100100},{9'b111111000},{9'b010101000},{9'b001000110},{9'b000100110},{9'b101010010},{9'b101011100},{9'b001010010},{9'b001001000},{9'b001010000},{9'b100100011},{9'b001010111},{9'b011101000},{9'b100100101},{9'b001000000},{9'b011100010},{9'b111100000},{9'b001000110},{9'b111001110},{9'b000100100},{9'b101001110},{9'b001000101},{9'b100011000},{9'b110110111},{9'b010000100},{9'b011110110},{9'b100001111},{9'b000001001},{9'b110010000},{9'b000011001},{9'b101111010},{9'b000110010},{9'b000011110},{9'b100000100},{9'b011011010},{9'b000110011},{9'b011010111},{9'b001000011},{9'b110100011},{9'b010111011},{9'b100110111},{9'b001101010},{9'b111010010},{9'b100110101},{9'b000101010},{9'b100001001},{9'b100111000},{9'b000110101},{9'b010001110},{9'b111101000},{9'b110110001},{9'b110000010},{9'b011100000},{9'b010001110},{9'b001011000},{9'b111101011},{9'b010010100},{9'b000111000},{9'b110101000},{9'b111010100},{9'b010001110},{9'b010001000},{9'b010011100},{9'b101001011},{9'b001011001},{9'b010100011},{9'b101111011},{9'b011110101},{9'b101100010},{9'b011101100},{9'b000100101},{9'b110001101},{9'b101011101},{9'b000101111},{9'b101111010},{9'b000110000},{9'b101010000},{9'b111001111},{9'b010000010},{9'b111000010},{9'b111100000},{9'b011000110},{9'b111100110},{9'b000010010},{9'b111110100},{9'b000100000},{9'b010001101},{9'b011101100},{9'b011010000},{9'b100110000},{9'b101101010},{9'b001111000},{9'b010100100},{9'b100111100},{9'b110110010},{9'b110110000},{9'b111110011},{9'b100101100},{9'b010101101},{9'b000010101},{9'b001100010},{9'b000010101},{9'b000011101},{9'b000001101},{9'b010101111},{9'b101111100},{9'b100011001},{9'b101100011},{9'b000100101},{9'b111000100},{9'b101110001},{9'b111110011},{9'b110011011},{9'b001101011},{9'b011001001},{9'b001010001},{9'b011110110},{9'b001010001},{9'b010101011},{9'b101011011},{9'b010010110},{9'b111111010},{9'b111001000},{9'b101110101},{9'b011011111},{9'b000001100},{9'b011000011},{9'b110111000},{9'b111110100},{9'b111010100},{9'b001111111},{9'b000100110},{9'b110001010},{9'b011011010},{9'b100111110},{9'b011101001},{9'b011111111},{9'b111110000},{9'b100000100},{9'b001110000},{9'b000100011},{9'b100101010},{9'b101101001},{9'b111110110},{9'b001011111},{9'b000000011},{9'b001100000},{9'b101101100},{9'b000100011},{9'b110101010},{9'b110000110},{9'b111001111},{9'b110001111},{9'b001101101},{9'b100001110},{9'b100110111},{9'b101000111},{9'b110100100},{9'b010000011},{9'b001000010},{9'b101110111},{9'b110000111},{9'b111000010},{9'b000110111},{9'b110101101},{9'b001100111},{9'b110110111},{9'b100011011},{9'b000110100},{9'b000010110},{9'b011101111},{9'b100100111},{9'b001100111},{9'b111101111},{9'b101010000},{9'b111001100},{9'b111010110},{9'b100101000},{9'b100110011},{9'b110010010},{9'b101101100},{9'b111011000},{9'b111011100},{9'b010010101},{9'b101011000},{9'b011010101},{9'b111100100},{9'b111001010},{9'b010000000},{9'b110001101},{9'b000110001},{9'b110001000},{9'b011001100},{9'b111001100},{9'b111111111},{9'b101011110},{9'b000110011},{9'b100011110},{9'b100100101},{9'b100001100},{9'b001111010},{9'b110001101},{9'b101101011},{9'b100100011},{9'b000010110},{9'b001101010},{9'b011001000},{9'b010000110},{9'b000001100},{9'b011111110},{9'b001100000},{9'b101100110},{9'b101111000},{9'b010001000},{9'b000110100},{9'b100101011},{9'b011001010},{9'b110001101},{9'b111100100},{9'b010001011},{9'b010101010},{9'b011011101},{9'b100100110},{9'b010000000},{9'b001010011},{9'b100010101},{9'b101111111},{9'b111010101},{9'b000010110},{9'b110110000},{9'b000000110},{9'b010110011},{9'b001100101},{9'b011101110},{9'b011001100},{9'b100101000},{9'b010001000},{9'b110000101},{9'b011111001},{9'b000010011},{9'b000001011},{9'b011110011},{9'b100000110},{9'b001111110},{9'b011010011},{9'b110101010},{9'b011101111},{9'b011101011},{9'b111101010},{9'b011011100},{9'b110000010},{9'b011010010},{9'b010001101},{9'b011111000},{9'b011100010},{9'b010111100},{9'b110010111},{9'b001011011},{9'b010110101},{9'b110011000},{9'b011000000},{9'b111111010},{9'b111100010},{9'b000100111},{9'b011110010},{9'b011110101},{9'b100010011},{9'b000001111},{9'b110111111},{9'b110001110},{9'b010001011},{9'b100010100},{9'b010011010},{9'b000010001},{9'b110001001},{9'b001110110},{9'b101111110},{9'b100001001},{9'b110011011},{9'b101100101},{9'b001001000},{9'b110101111},{9'b101001100},{9'b011010100},{9'b011000100},{9'b110011110},{9'b010010011},{9'b101100110},{9'b011010101},{9'b011000010},{9'b100011010},{9'b000100010},{9'b011001111},{9'b101101010},{9'b111110001},{9'b101101011},{9'b111110001},{9'b000000001},{9'b001010100},{9'b010001010},{9'b100110110},{9'b111011011},{9'b111110011},{9'b010101000},{9'b000001011},{9'b011110111},{9'b110011110},{9'b100101100},{9'b001010011},{9'b000101100},{9'b001100111},{9'b101101100},{9'b001110010},{9'b001000110},{9'b010110110},{9'b001001000},{9'b001010000},{9'b011001000},{9'b110100010},{9'b110111100},{9'b110001111},{9'b101011100},{9'b111111101},{9'b110111011},{9'b100011000},{9'b101111101},{9'b000011110},{9'b101010011},{9'b100001100},{9'b100110010},{9'b010101100},{9'b110010000},{9'b011101100},{9'b111111001},{9'b000111011},{9'b001110110},{9'b001101010},{9'b010000001},{9'b101101111},{9'b011011111},{9'b001000011},{9'b001111000},{9'b011000010},{9'b100001011},{9'b000101011},{9'b111001100},{9'b010110001},{9'b100111100},{9'b001000100},{9'b110011110},{9'b010011110},{9'b101100110},{9'b011010101},{9'b111000011},{9'b100111101},{9'b110110101},{9'b011010111},{9'b000000011},{9'b100000001},{9'b011100010},{9'b000101110},{9'b101111001},{9'b101011000},{9'b100001011},{9'b100011000},{9'b010010001},{9'b100000111},{9'b000110001},{9'b001100101},{9'b001101111},{9'b010100101},{9'b110010000},{9'b101100111},{9'b111100010},{9'b110001011},{9'b010000010},{9'b100000100},{9'b110111001},{9'b110001101},{9'b101001010},{9'b110001010},{9'b101010110},{9'b110100011},{9'b111100101},{9'b000101110},{9'b111111101},{9'b100100001},{9'b000000110},{9'b110111001},{9'b011110001},{9'b011110001},{9'b000110101},{9'b011111001},{9'b011100001},{9'b100110010},{9'b011110111},{9'b010011101},{9'b000100110},{9'b001000010},{9'b001100010},{9'b100101100},{9'b001111001},{9'b101000110},{9'b001000101},{9'b111000100},{9'b101000000},{9'b001011000},{9'b100010000},{9'b110011000},{9'b010100010},{9'b101001010},{9'b110110110},{9'b101011111},{9'b011011100},{9'b100000010},{9'b100101010},{9'b010111100},{9'b001000110},{9'b110110010},{9'b111010000},{9'b001000100},{9'b010010000},{9'b000011000},{9'b000111011},{9'b011000000},{9'b110001110},{9'b101111110},{9'b011011111},{9'b110001110},{9'b110110111},{9'b011010110},{9'b010001110},{9'b011100001},{9'b000000100},{9'b010100100},{9'b001010011},{9'b000111000},{9'b011100110},{9'b000101001},{9'b101010010},{9'b101101110},{9'b101000010},{9'b101101000},{9'b001000000},{9'b000010101},{9'b100111000},{9'b110100101},{9'b100000001},{9'b001010011},{9'b110001011},{9'b100001011},{9'b110010100},{9'b101110001},{9'b010111000},{9'b001000100},{9'b111001100},{9'b011001101},{9'b111100111},{9'b111011100},{9'b010100100},{9'b101101100},{9'b000101001},{9'b010000110},{9'b111100100},{9'b100110101},{9'b101010110},{9'b100001011},{9'b010100001},{9'b101110011},{9'b011100110},{9'b011101001},{9'b001011111},{9'b011110100},{9'b101101101},{9'b000001101},{9'b100010010},{9'b010110111},{9'b101001000},{9'b101111010},{9'b001111011},{9'b001000010},{9'b000101101},{9'b001000100},{9'b010111001},{9'b111001011},{9'b011111001},{9'b010110101},{9'b011110011},{9'b000010001},{9'b011111101},{9'b110100011},{9'b000001000},{9'b001011010},{9'b000011000},{9'b001000100},{9'b110100001},{9'b011001010},{9'b000110100},{9'b011110101},{9'b010101011},{9'b000111011},{9'b011100011},{9'b010000101},{9'b111110111},{9'b000001000},{9'b110000000},{9'b100110110},{9'b101100111},{9'b100100100},{9'b000101010},{9'b010111001},{9'b010001100},{9'b110010000},{9'b110000000},{9'b110100000},{9'b011000010},{9'b000111101},{9'b101001111},{9'b101001110},{9'b011001000},{9'b001100110},{9'b000011001},{9'b011000001},{9'b010011010},{9'b110110001},{9'b010111011},{9'b100001111},{9'b010010001},{9'b000001011},{9'b000011001},{9'b110010101},{9'b101011001},{9'b101100011},{9'b011101000},{9'b010010111},{9'b011001110},{9'b001100100},{9'b100101001},{9'b000101000},{9'b010001000},{9'b101110011},{9'b011010100},{9'b011010100},{9'b101101111},{9'b110111100},{9'b010111010},{9'b011010000},{9'b010101010},{9'b000110100},{9'b010110011},{9'b010000010},{9'b000101001},{9'b110011000},{9'b100001000},{9'b101011001},{9'b110111100},{9'b101000101},{9'b001111100},{9'b111001110},{9'b101111010},{9'b101110110},{9'b000010000},{9'b101000110},{9'b000101100},{9'b011000111},{9'b101000111},{9'b011001101},{9'b101100101},{9'b001010010},{9'b001110110},{9'b101101101},{9'b110001101},{9'b000110001},{9'b101011010},{9'b100111010},{9'b000100100},{9'b011001011},{9'b000010001},{9'b110010111},{9'b000011010},{9'b110110100},{9'b001011100},{9'b000010010},{9'b100111010},{9'b111001010},{9'b111011111},{9'b110101100},{9'b111000100},{9'b001110000},{9'b000100010},{9'b111001111},{9'b001111100},{9'b101001111},{9'b111101011},{9'b000000101},{9'b011111010},{9'b001010101},{9'b001000001},{9'b001010110},{9'b101111010},{9'b010100011},{9'b010110001},{9'b100010010},{9'b111011111},{9'b001001010},{9'b000100001},{9'b101010000},{9'b100011010},{9'b010100001},{9'b001100111},{9'b100110000},{9'b001001010},{9'b000001100},{9'b010111101},{9'b000101100},{9'b000000001},{9'b011010110},{9'b001101011},{9'b001010111},{9'b110100111},{9'b001100101},{9'b101001010},{9'b101101110},{9'b010011011},{9'b101000010},{9'b011111010},{9'b101101001},{9'b011100000},{9'b011111111},{9'b011001100},{9'b001000011},{9'b000110101},{9'b010011000},{9'b011111110},{9'b110000000},{9'b011111011},{9'b001000111},{9'b001101110},{9'b110011110},{9'b000111011},{9'b100111010},{9'b110110100},{9'b111111011},{9'b010101101},{9'b101101010},{9'b011100111},{9'b111000110},{9'b110110000},{9'b111001100},{9'b101111000},{9'b110110000},{9'b111010101},{9'b011100101},{9'b010110001},{9'b100101011},{9'b010111001},{9'b110101011},{9'b111111011},{9'b101100101},{9'b011010110},{9'b001010000},{9'b000111000},{9'b001000110},{9'b100000110},{9'b000111110},{9'b001100001},{9'b011100010},{9'b110111000},{9'b010110110},{9'b100000001},{9'b000110111},{9'b000010010},{9'b001110101},{9'b011011100},{9'b100100100},{9'b111001000},{9'b100101100},{9'b110111101},{9'b010111111},{9'b110100101},{9'b001011000},{9'b110001110},{9'b011110110},{9'b011000100},{9'b111010011},{9'b110100110},{9'b111000110},{9'b000001101},{9'b011001001},{9'b001110011},{9'b000000100},{9'b001101001},{9'b011010011},{9'b001100011},{9'b001011111},{9'b101111001},{9'b100110101},{9'b110110001},{9'b101110011},{9'b110110101},{9'b101100000},{9'b001010001},{9'b110010010},{9'b100111100},{9'b100010010},{9'b111001011},{9'b011101101},{9'b010111010},{9'b110000101},{9'b011001000},{9'b001000101},{9'b110001110},{9'b010011101},{9'b011001101},{9'b001010010},{9'b000000100},{9'b111010011},{9'b111011001},{9'b010011010},{9'b111000010},{9'b010011001},{9'b111011010},{9'b011111110},{9'b100100000},{9'b010110001},{9'b100100100},{9'b000001011},{9'b010010101},{9'b010010110},{9'b000110010},{9'b111110110},{9'b001110000},{9'b110010001},{9'b001011100},{9'b011111010},{9'b000101011},{9'b101011001},{9'b010101101},{9'b011011011},{9'b011101010},{9'b010100101},{9'b000000011},{9'b100000111},{9'b000110000},{9'b101010100},{9'b010111101},{9'b100111101},{9'b011010011},{9'b001011101},{9'b110001100},{9'b100111101},{9'b011111011},{9'b101110111},{9'b100111110},{9'b010110111},{9'b101010000},{9'b011100001},{9'b110011011},{9'b101010111},{9'b110101001},{9'b100110101},{9'b000110101},{9'b101111001},{9'b110111111},{9'b101101001},{9'b001000001},{9'b000010000},{9'b010101011},{9'b100010000},{9'b100101010},{9'b010101010},{9'b010001100},{9'b010101101},{9'b010110101},{9'b011101111},{9'b010101001},{9'b001011101},{9'b101001101},{9'b111011011},{9'b100001000},{9'b000100100},{9'b100110010},{9'b010101000},{9'b000001100},{9'b110100001},{9'b100000110},{9'b001110001},{9'b110011111},{9'b111110001},{9'b100101011},{9'b011110001},{9'b011100101},{9'b101111111},{9'b001011111},{9'b100010010},{9'b001011001},{9'b010001011},{9'b010000111},{9'b011001011},{9'b010010011},{9'b100011000},{9'b011011001},{9'b010111001},{9'b001010011},{9'b001111010},{9'b010010001},{9'b001011010},{9'b110010111},{9'b110101110},{9'b011000011},{9'b000110010},{9'b100001110},{9'b010001000},{9'b101101010},{9'b010001100},{9'b011111000},{9'b101011100},{9'b000001111},{9'b001010101},{9'b011001001},{9'b011110011},{9'b001111010},{9'b000000111},{9'b001110111},{9'b110101100},{9'b100001000},{9'b100001000},{9'b101101001},{9'b011110101},{9'b100100101},{9'b000111111},{9'b001100011},{9'b001111011},{9'b000101111},{9'b001101110},{9'b101111101},{9'b101001010},{9'b010001001},{9'b100000010},{9'b010001101},{9'b011000101},{9'b011010010},{9'b111001101},{9'b011001110},{9'b101001101},{9'b001001000},{9'b111101011},{9'b101110100},{9'b001011010},{9'b100001101},{9'b011011010},{9'b110111000},{9'b010100111},{9'b110111011},{9'b011010000},{9'b000110111},{9'b111111100},{9'b110000101},{9'b100101111},{9'b011110110},{9'b010000100},{9'b101010001},{9'b100111110},{9'b011100000},{9'b100100111},{9'b111011100},{9'b101100101},{9'b000000100},{9'b101001001},{9'b101001111},{9'b111100000},{9'b100001010},{9'b010011011},{9'b110110110},{9'b111110111},{9'b011010100},{9'b111001111},{9'b111111001},{9'b100100001},{9'b100010111},{9'b010011010},{9'b100010100},{9'b110111101},{9'b110011010},{9'b110101001},{9'b011101101},{9'b101110101},{9'b100010001},{9'b100000011},{9'b111000010},{9'b101010001},{9'b001001001},{9'b111110101},{9'b110010111},{9'b110111111},{9'b111100101},{9'b011111110},{9'b101011001},{9'b111100011},{9'b000000001},{9'b001110110},{9'b111010001},{9'b000001111},{9'b111011000},{9'b100100101},{9'b100011010},{9'b001010101},{9'b111100010},{9'b101001011},{9'b111000000},{9'b111011010},{9'b010101011},{9'b100001110},{9'b001111000},{9'b010100101},{9'b010110001},{9'b010100101},{9'b101101101},{9'b001011000},{9'b010000100},{9'b000111101},{9'b010011000},{9'b011110000},{9'b100010001},{9'b101011101},{9'b100001010},{9'b110011001},{9'b111111111},{9'b010010000},{9'b000110101},{9'b001110001},{9'b111011101},{9'b110011010},{9'b010111001},{9'b100000101},{9'b010010110},{9'b100010110},{9'b100000010},{9'b000010110},{9'b001101010},{9'b100110001},{9'b111000011},{9'b110100000},{9'b000001000},{9'b101011101},{9'b111110101},{9'b111101010},{9'b101100111},{9'b100010100},{9'b000100101},{9'b111111001},{9'b101001110},{9'b001111011},{9'b001010010},{9'b010010110},{9'b001000000},{9'b101110110},{9'b100101110},{9'b110000110},{9'b000111101},{9'b010110011},{9'b101011001},{9'b100111101},{9'b010101001},{9'b011110110},{9'b011010011},{9'b110111110},{9'b101100101},{9'b011101110},{9'b010111011},{9'b100001101},{9'b100111010},{9'b001100101},{9'b111111101},{9'b000110111},{9'b101110111},{9'b001111111},{9'b110000000},{9'b100011111},{9'b001100010},{9'b101011000},{9'b100011001},{9'b100111110},{9'b100111111},{9'b011011110},{9'b110011010},{9'b101000100},{9'b000010001},{9'b101011101},{9'b101101010},{9'b010000101},{9'b101101110},{9'b110000010},{9'b000011001},{9'b100010001},{9'b010000001},{9'b101010111},{9'b001100001},{9'b011001101},{9'b111101100},{9'b100010010},{9'b000010100},{9'b111010111},{9'b011010111},{9'b000000101},{9'b110110111},{9'b001001101},{9'b100000101},{9'b000100001},{9'b010000100},{9'b011000100},{9'b010101100},{9'b010000011},{9'b011110111},{9'b000001110},{9'b101001100},{9'b111111101},{9'b100110101},{9'b010110111},{9'b111101111},{9'b101010010},{9'b111101111},{9'b100101010},{9'b100010101},{9'b001101001},{9'b011001001},{9'b100100001},{9'b111101011},{9'b111010110},{9'b110101011},{9'b101111110},{9'b101111101},{9'b010101100},{9'b111101011},{9'b100000100},{9'b101111111},{9'b001100011},{9'b110100001},{9'b010111010},{9'b110010011},{9'b101001001},{9'b111111010},{9'b011111100},{9'b111010110},{9'b110000000},{9'b000000101},{9'b100010100},{9'b110001101},{9'b010010110},{9'b010010010},{9'b101000011},{9'b100110000},{9'b001100110},{9'b110101101},{9'b010100010},{9'b100110111},{9'b101111101},{9'b001011110},{9'b101101100},{9'b000011110},{9'b010100001},{9'b111111110},{9'b010111001},{9'b100001100},{9'b000111000},{9'b100111000},{9'b011111110},{9'b111000101},{9'b011011111},{9'b111110010},{9'b101000011},{9'b011100111},{9'b011011101},{9'b110000001},{9'b000100010},{9'b001000011},{9'b101111100},{9'b001000110},{9'b111110110},{9'b101100001},{9'b110010011},{9'b001101100},{9'b101111010},{9'b110100110},{9'b000001100},{9'b000010111},{9'b011001011},{9'b100111010},{9'b001000011},{9'b010100011},{9'b001010111},{9'b000011100},{9'b110100010},{9'b001111010},{9'b100110010},{9'b010011011},{9'b000001110},{9'b110111110},{9'b101011000},{9'b101110111},{9'b010100110},{9'b011110100},{9'b101000101},{9'b100000111},{9'b111111110},{9'b110000001},{9'b001001010},{9'b111010101},{9'b010110111},{9'b111011000},{9'b111011110},{9'b111010111},{9'b110101011},{9'b010010110},{9'b001011110},{9'b100101101},{9'b000101011},{9'b110100101},{9'b000111001},{9'b000000010},{9'b000010001},{9'b111011000},{9'b110111100},{9'b000010101},{9'b100010000},{9'b100111100},{9'b111110000},{9'b100001100},{9'b000011000},{9'b100100101},{9'b101011100},{9'b110111001},{9'b110000101},{9'b101011100},{9'b101111011},{9'b101000011},{9'b101001011},{9'b010001100},{9'b000101101},{9'b010010101},{9'b101001010},{9'b110011010},{9'b011100011},{9'b011000001},{9'b101100010},{9'b110010011},{9'b011100010},{9'b111001101},{9'b001011101},{9'b000100101},{9'b101101100},{9'b111000010},{9'b110110000},{9'b101011100},{9'b111111010},{9'b010100101},{9'b001001101},{9'b110001001},{9'b001110101},{9'b100011011},{9'b101111011},{9'b010101111},{9'b011011111},{9'b010110000},{9'b111111001},{9'b000010001},{9'b100001111},{9'b000110101},{9'b001100110},{9'b100111101},{9'b110110011},{9'b000110011},{9'b011110110},{9'b010001010},{9'b011110000},{9'b011001000},{9'b011110011},{9'b100101100},{9'b011000110},{9'b000101110},{9'b101100010},{9'b110110111},{9'b010111101},{9'b011110010},{9'b111010100},{9'b000001111},{9'b000000011},{9'b010111000},{9'b101110001},{9'b100100011},{9'b110111100},{9'b011000011},{9'b000011111},{9'b011011100},{9'b100010000},{9'b000110000},{9'b100101011},{9'b010111110},{9'b011100110},{9'b100000101},{9'b111101011},{9'b010010000},{9'b110001000},{9'b001100101},{9'b111111100},{9'b001100001},{9'b010000010},{9'b101100111},{9'b001001000},{9'b010000110},{9'b000001010},{9'b000101000},{9'b000100011},{9'b101101001},{9'b100100101},{9'b111001010},{9'b100111110},{9'b111111100},{9'b011111010},{9'b011000110},{9'b000001111},{9'b111001010},{9'b100100010},{9'b100010110},{9'b101101010},{9'b011110111},{9'b000110101},{9'b101101110},{9'b001110011},{9'b001110010},{9'b011001101},{9'b100011101},{9'b011011110},{9'b101100001},{9'b100001100},{9'b011111000},{9'b001000000},{9'b111100101},{9'b101111111},{9'b010110101},{9'b010101101},{9'b111101001},{9'b101011100},{9'b100111110},{9'b100010001},{9'b001010010},{9'b101100110},{9'b001111000},{9'b110010110},{9'b001110111},{9'b110101111},{9'b100110110},{9'b011010001},{9'b100011110},{9'b101111001},{9'b011101000},{9'b110110101},{9'b111011110},{9'b111001011},{9'b000011110},{9'b101011001},{9'b010111110},{9'b011100100},{9'b100011001},{9'b010100000},{9'b101101100},{9'b010010100},{9'b110101110},{9'b001011100},{9'b010000000},{9'b010100100},{9'b001001110},{9'b000001000},{9'b001011110},{9'b100001011},{9'b010101100},{9'b011110110},{9'b110111001},{9'b011011010},{9'b100110101},{9'b010001011},{9'b010100011},{9'b110110110},{9'b100001000},{9'b100011010},{9'b110010110},{9'b001110110},{9'b010111010},{9'b000100111},{9'b100010000},{9'b100010000},{9'b110101011},{9'b010000000},{9'b011111010},{9'b111011101},{9'b101001001},{9'b000011111},{9'b111100011},{9'b001011000},{9'b001111110},{9'b000101110},{9'b010100100},{9'b110010011},{9'b100101101},{9'b110001010},{9'b101111101},{9'b100101001},{9'b001011100},{9'b001001101},{9'b011000010},{9'b010010011},{9'b001100000},{9'b011001010},{9'b001000100},{9'b100111001},{9'b110011011},{9'b100110001},{9'b101110011},{9'b101011000},{9'b111011111},{9'b000100010},{9'b100110101},{9'b110101000},{9'b101101101},{9'b001111110},{9'b101110100},{9'b110101010},{9'b111110010},{9'b001110110},{9'b001001101},{9'b111001010},{9'b011011100},{9'b011001111},{9'b011010010},{9'b110101010},{9'b100110101},{9'b101111100},{9'b010001110},{9'b110010110},{9'b011101111},{9'b000110111},{9'b101101001},{9'b111111001},{9'b110000001},{9'b110100000},{9'b010000011},{9'b001100010},{9'b011100000},{9'b100010010},{9'b101110110},{9'b110010000},{9'b111111001},{9'b110010000},{9'b101001010},{9'b110011010},{9'b011110001},{9'b001001100},{9'b011110000},{9'b110100011},{9'b000101101},{9'b001100110},{9'b101000111},{9'b101000000},{9'b011011011},{9'b000111010},{9'b010010000},{9'b111010100},{9'b101000110},{9'b010001001},{9'b110110110},{9'b010100100},{9'b100101000},{9'b001001110},{9'b110010010},{9'b001000100},{9'b000111101},{9'b010010000},{9'b001111011},{9'b111101110},{9'b100101100},{9'b101100010},{9'b011001101},{9'b110111110},{9'b001100000},{9'b000011000},{9'b010011010},{9'b010010100},{9'b010100000},{9'b110110000},{9'b111110100},{9'b011110101},{9'b100001101},{9'b100001001},{9'b100011101},{9'b000110101},{9'b100011101},{9'b010101001},{9'b110111001},{9'b001110111},{9'b010101110},{9'b001100101},{9'b001110101},{9'b001110100},{9'b011101011},{9'b001111001},{9'b111000111},{9'b010110000},{9'b011010010},{9'b000001101},{9'b100100011},{9'b011001100},{9'b110011101},{9'b100011001},{9'b110111001},{9'b101011101},{9'b010001011},{9'b100011011},{9'b000101111},{9'b010001111},{9'b010110000},{9'b100110000},{9'b111001111},{9'b101001001},{9'b111001001},{9'b110011111},{9'b001000111},{9'b100101000},{9'b001111000},{9'b111101111},{9'b001100011},{9'b010101110},{9'b101110110},{9'b101100111},{9'b001011100},{9'b110011010},{9'b101010010},{9'b110110110},{9'b101100100},{9'b000100111},{9'b011000010},{9'b101101010},{9'b111001000},{9'b100011010},{9'b100111100},{9'b001100111},{9'b101001111},{9'b110110010},{9'b001100000},{9'b100100001},{9'b010000011},{9'b001111100},{9'b001101011},{9'b001001111},{9'b001010111},{9'b111011100},{9'b011101110},{9'b101111110},{9'b110001111},{9'b001011000},{9'b001010001},{9'b011111100},{9'b101011000},{9'b110000010},{9'b000100010},{9'b110101111},{9'b100011010},{9'b110010100},{9'b101010000},{9'b111001111},{9'b110110011},{9'b111010111},{9'b000111011},{9'b100110011},{9'b100111010},{9'b011111010},{9'b110111110},{9'b111101111},{9'b001001000},{9'b001000100},{9'b001110010},{9'b101010001},{9'b100110000},{9'b111001000},{9'b011010001},{9'b110001111},{9'b111100110},{9'b111001100},{9'b111001110},{9'b111010101},{9'b011101111},{9'b001011000},{9'b110011110},{9'b001001011},{9'b010111010},{9'b101001000},{9'b011101010},{9'b011011111},{9'b000101000},{9'b011011100},{9'b001000100},{9'b111110110},{9'b011110100},{9'b010100010},{9'b111000110},{9'b101111001},{9'b111111010},{9'b110111000},{9'b001000110},{9'b000100100},{9'b010001011},{9'b001110010},{9'b110101011},{9'b100111000},{9'b100101111},{9'b111101101},{9'b111101111},{9'b010111101},{9'b100011101},{9'b101001110},{9'b011111110},{9'b101010001},{9'b011101010},{9'b001011101},{9'b011010001},{9'b101111010},{9'b111111000},{9'b010000010},{9'b110001111},{9'b011101011},{9'b001001011},{9'b011101111},{9'b101011101},{9'b001001010},{9'b110111000},{9'b101001110},{9'b101110000},{9'b001010110},{9'b011111100},{9'b101111111},{9'b101110010},{9'b011100000},{9'b010011011},{9'b100011100},{9'b100001101},{9'b110011000},{9'b111101010},{9'b010001100},{9'b011110111},{9'b001101101},{9'b000111101},{9'b000110011},{9'b000100000},{9'b011101100},{9'b000110011},{9'b100001100},{9'b101110110},{9'b111000010},{9'b000011011},{9'b110110110},{9'b100101010},{9'b001110110},{9'b110001100},{9'b110010010},{9'b001101111},{9'b110100011},{9'b011110101},{9'b101110100},{9'b010010010},{9'b100101111},{9'b111001110},{9'b110001100},{9'b000101111},{9'b011100100},{9'b100001001},{9'b101011111},{9'b100011110},{9'b010101010},{9'b010111001},{9'b110001010},{9'b111000100},{9'b111001111},{9'b010101010},{9'b100001011},{9'b101010001},{9'b001100100},{9'b100001000},{9'b110110101},{9'b110010000},{9'b001111010},{9'b111001111},{9'b001000110},{9'b110010101},{9'b001100110},{9'b011011100},{9'b001101001},{9'b011001011},{9'b011111111},{9'b111110000},{9'b111001110},{9'b100010011},{9'b100001111},{9'b000011110},{9'b001000001},{9'b111111101},{9'b110000011},{9'b010001100},{9'b010100011},{9'b010100011},{9'b001101010},{9'b000111101},{9'b101110011},{9'b000101010},{9'b110011101},{9'b110111100},{9'b101001111},{9'b010111001},{9'b101010111},{9'b101001110},{9'b011011101},{9'b011010010},{9'b000111101},{9'b110011101},{9'b100011000},{9'b100000101},{9'b010001100},{9'b011010010},{9'b101110100},{9'b011000011},{9'b001110001},{9'b100110011},{9'b111111101},{9'b010011001},{9'b110010110},{9'b001101001},{9'b010100111},{9'b100111011},{9'b011011000},{9'b010110010},{9'b000001011},{9'b110011100},{9'b111111001},{9'b010010000},{9'b010011100},{9'b011101110},{9'b101110110},{9'b011110110},{9'b111110111},{9'b100101010},{9'b000011000},{9'b111110100},{9'b101111110},{9'b011110111},{9'b101010110},{9'b001100001},{9'b111111001},{9'b110101100},{9'b011110000},{9'b110110101},{9'b000100011},{9'b110101001},{9'b000110000},{9'b111101000},{9'b110110010},{9'b101111110},{9'b010011010},{9'b001011000},{9'b011010101},{9'b010001010},{9'b011111100},{9'b010101100},{9'b100110011},{9'b000010010},{9'b001101010},{9'b000010101},{9'b110101011},{9'b001111010},{9'b100011110},{9'b000110011},{9'b101110011},{9'b000110010},{9'b110011010},{9'b101111010},{9'b111100111},{9'b011101011},{9'b000000110},{9'b100001011},{9'b110011110},{9'b100001010},{9'b111101110},{9'b110011100},{9'b010011010},{9'b100111000},{9'b001100110},{9'b110101010},{9'b111110110},{9'b101011111},{9'b001111001},{9'b001110111},{9'b000100110},{9'b100101100},{9'b110011001},{9'b011101110},{9'b111001100},{9'b111101011},{9'b000010110},{9'b001111000},{9'b100011101},{9'b100011000},{9'b111010001},{9'b000101111},{9'b111001011},{9'b011011010},{9'b010011000},{9'b011101110},{9'b001100110},{9'b011001111},{9'b101010011},{9'b011110011},{9'b110101001},{9'b101111110},{9'b000110100},{9'b011111010},{9'b101110111},{9'b010101010},{9'b101001011},{9'b110001110},{9'b111111001},{9'b011011101},{9'b010101100},{9'b001001000},{9'b101110110},{9'b111111001},{9'b010011110},{9'b111101111},{9'b010000110},{9'b100101001},{9'b100101000},{9'b010111011},{9'b110111000},{9'b001101001},{9'b000010111},{9'b110111101},{9'b110110111},{9'b100000000},{9'b100001110},{9'b011111000},{9'b001000100},{9'b101011110},{9'b010010010},{9'b010010011},{9'b101110101},{9'b110011011},{9'b110100011},{9'b110101100},{9'b001110101},{9'b011001101},{9'b010101001},{9'b100101101},{9'b000111010},{9'b010000011},{9'b100000111},{9'b011011000}};
assign weight_o_2 = {{9'b010100011},{9'b001100111},{9'b111000000},{9'b110100001},{9'b011100001},{9'b001101001},{9'b011100010},{9'b100011000},{9'b000111011},{9'b110001101},{9'b101101111},{9'b111011100},{9'b100000010},{9'b011001011},{9'b001001111},{9'b100000101},{9'b110010101},{9'b001110011},{9'b000011110},{9'b000110010},{9'b000001000},{9'b100110111},{9'b101011110},{9'b000100001},{9'b000010100},{9'b100101001},{9'b001010011},{9'b111001100},{9'b010101011},{9'b110001111},{9'b011110100},{9'b100011000},{9'b011111100},{9'b001101000},{9'b010100111},{9'b010101000},{9'b010001111},{9'b100101000},{9'b111000100},{9'b010010110},{9'b100100100},{9'b000110011},{9'b101111100},{9'b000011111},{9'b110101010},{9'b111010100},{9'b100011011},{9'b110110101},{9'b110010000},{9'b100010100},{9'b011110010},{9'b110010110},{9'b001001011},{9'b111011110},{9'b111011010},{9'b111100110},{9'b100001001},{9'b111110011},{9'b111001101},{9'b000010001},{9'b100011101},{9'b011010011},{9'b100000101},{9'b110101110},{9'b011110100},{9'b010010100},{9'b100000100},{9'b011010000},{9'b001101110},{9'b110110011},{9'b000100111},{9'b111111110},{9'b001001100},{9'b011000110},{9'b110011100},{9'b011100011},{9'b101000001},{9'b111101110},{9'b101111011},{9'b101000100},{9'b011001011},{9'b011100111},{9'b011011001},{9'b101101110},{9'b011011010},{9'b010010001},{9'b111100011},{9'b100001000},{9'b110011111},{9'b010111111},{9'b100101111},{9'b011100011},{9'b001010011},{9'b111000110},{9'b011010100},{9'b100011000},{9'b001010101},{9'b111110110},{9'b110101110},{9'b011001010},{9'b000111110},{9'b100001111},{9'b101000110},{9'b110111011},{9'b101000100},{9'b100111001},{9'b100101100},{9'b110011111},{9'b010110010},{9'b100000111},{9'b010011010},{9'b111100001},{9'b100010100},{9'b100010110},{9'b101100010},{9'b011110111},{9'b010110011},{9'b111100101},{9'b101001111},{9'b000010111},{9'b010010100},{9'b001100000},{9'b011001111},{9'b010010011},{9'b000000101},{9'b010010011},{9'b010011010},{9'b111001100},{9'b000010101},{9'b000111000},{9'b000011110},{9'b001110000},{9'b101101000},{9'b110110110},{9'b100001100},{9'b110011001},{9'b100011011},{9'b100101000},{9'b001000001},{9'b110011111},{9'b000111010},{9'b000111001},{9'b010010111},{9'b010000000},{9'b101100001},{9'b101000011},{9'b001010101},{9'b101101110},{9'b011101000},{9'b111111010},{9'b001011110},{9'b000101001},{9'b100111010},{9'b000101000},{9'b000110000},{9'b010100000},{9'b100111011},{9'b111000011},{9'b011000000},{9'b000110010},{9'b001111100},{9'b110110100},{9'b111011100},{9'b110001010},{9'b000011111},{9'b000000110},{9'b101101111},{9'b100000011},{9'b010101100},{9'b000111000},{9'b001011110},{9'b111100000},{9'b101110010},{9'b001000110},{9'b011000111},{9'b001110010},{9'b101101110},{9'b010111010},{9'b110110110},{9'b000110100},{9'b110100111},{9'b011110110},{9'b100011000},{9'b111100110},{9'b100010100},{9'b100111101},{9'b000011010},{9'b010010000},{9'b101011111},{9'b111001101},{9'b001110111},{9'b000000010},{9'b010111000},{9'b001111011},{9'b111001000},{9'b010101001},{9'b011000001},{9'b111001100},{9'b011010111},{9'b110100001},{9'b011101100},{9'b101101111},{9'b001101000},{9'b110011010},{9'b011001001},{9'b100011101},{9'b110111111},{9'b011000110},{9'b011000001},{9'b101111111},{9'b111010101},{9'b101001100},{9'b011000100},{9'b111011010},{9'b111111101},{9'b001101001},{9'b100011101},{9'b011101111},{9'b100100110},{9'b010001100},{9'b001101100},{9'b010111110},{9'b000110100},{9'b100011101},{9'b001110110},{9'b100011111},{9'b001010110},{9'b000111000},{9'b110011110},{9'b100110111},{9'b100010100},{9'b100100111},{9'b000101111},{9'b001010001},{9'b100111110},{9'b011010011},{9'b100110110},{9'b110000110},{9'b000011001},{9'b101001001},{9'b100100101},{9'b110010011},{9'b111100000},{9'b010101000},{9'b101001001},{9'b101000101},{9'b110011111},{9'b001101111},{9'b101111110},{9'b101111000},{9'b101000111},{9'b010011000},{9'b100111011},{9'b110011011},{9'b101011111},{9'b011101011},{9'b010111101},{9'b000111010},{9'b100011001},{9'b110011101},{9'b111000010},{9'b110011001},{9'b111010111},{9'b001101111},{9'b000010110},{9'b100000011},{9'b001111111},{9'b011101011},{9'b010011000},{9'b110001001},{9'b111110111},{9'b110101011},{9'b101000010},{9'b011101010},{9'b110110010},{9'b001110110},{9'b100111010},{9'b011010111},{9'b001101110},{9'b111011000},{9'b100110100},{9'b100111110},{9'b000001110},{9'b101101000},{9'b010000001},{9'b100001111},{9'b000011011},{9'b110111001},{9'b100101100},{9'b001111000},{9'b000110001},{9'b011010110},{9'b100111111},{9'b000101000},{9'b011000111},{9'b100111010},{9'b100011001},{9'b100110001},{9'b000011101},{9'b000010111},{9'b010001101},{9'b110110001},{9'b010001000},{9'b110000010},{9'b010011100},{9'b100011101},{9'b001010110},{9'b011110000},{9'b001001101},{9'b100111011},{9'b010111000},{9'b010011010},{9'b001000100},{9'b000000111},{9'b010101110},{9'b010100000},{9'b000000011},{9'b111111001},{9'b011100111},{9'b001100101},{9'b000101111},{9'b111100111},{9'b110001000},{9'b010100111},{9'b001011001},{9'b111110010},{9'b010100011},{9'b111110110},{9'b110000100},{9'b010000000},{9'b010010001},{9'b010100011},{9'b101011111},{9'b111100100},{9'b100000111},{9'b001001010},{9'b010010001},{9'b101101011},{9'b001010101},{9'b101101110},{9'b011000000},{9'b110111011},{9'b101100111},{9'b111000100},{9'b100110011},{9'b000101000},{9'b110110111},{9'b110101010},{9'b101000010},{9'b001111111},{9'b011100111},{9'b000010000},{9'b011110001},{9'b110110000},{9'b100001110},{9'b001011111},{9'b101110001},{9'b101101010},{9'b010011001},{9'b010101110},{9'b011010011},{9'b001100111},{9'b010010110},{9'b100111100},{9'b100111101},{9'b001001110},{9'b100010101},{9'b011101001},{9'b111010001},{9'b100000000},{9'b010000001},{9'b101101111},{9'b101011001},{9'b100010110},{9'b111100101},{9'b000010011},{9'b011001011},{9'b110011000},{9'b001010001},{9'b000011101},{9'b011110000},{9'b010000101},{9'b100011101},{9'b100111011},{9'b111111100},{9'b000101000},{9'b101101100},{9'b110011101},{9'b001001110},{9'b110010011},{9'b111001101},{9'b010011001},{9'b111101111},{9'b101011001},{9'b101111010},{9'b101101110},{9'b010100100},{9'b100010001},{9'b110001011},{9'b001001101},{9'b111000001},{9'b111101011},{9'b001011011},{9'b110101010},{9'b010010111},{9'b110100011},{9'b110000110},{9'b110001110},{9'b001100000},{9'b011010001},{9'b011001001},{9'b100011111},{9'b110000110},{9'b111111000},{9'b100110111},{9'b111000111},{9'b101100011},{9'b000111001},{9'b001110110},{9'b110011000},{9'b100111010},{9'b101010101},{9'b101111101},{9'b101110111},{9'b001010011},{9'b000101101},{9'b100101011},{9'b101111100},{9'b101010001},{9'b001000100},{9'b100011101},{9'b011100101},{9'b111010111},{9'b100000001},{9'b111110000},{9'b111111010},{9'b000110011},{9'b000111110},{9'b110101111},{9'b000101011},{9'b111110100},{9'b011011110},{9'b110010010},{9'b100101100},{9'b011110111},{9'b010101001},{9'b000110111},{9'b100000001},{9'b011111110},{9'b111100110},{9'b100001000},{9'b110101111},{9'b101101001},{9'b001110110},{9'b001100011},{9'b000111101},{9'b000011011},{9'b011100000},{9'b111110110},{9'b110001011},{9'b011000101},{9'b111010001},{9'b101000111},{9'b111011000},{9'b000000011},{9'b100010000},{9'b100011011},{9'b000101011},{9'b001100101},{9'b101111111},{9'b100101110},{9'b001111010},{9'b010010010},{9'b001001011},{9'b110111001},{9'b101100100},{9'b111010100},{9'b011101001},{9'b000011100},{9'b110010101},{9'b000101000},{9'b011011010},{9'b011001110},{9'b111011001},{9'b100001101},{9'b100111010},{9'b000000100},{9'b000001111},{9'b010110110},{9'b011011011},{9'b001011000},{9'b001000101},{9'b101010001},{9'b101000101},{9'b000000110},{9'b001010110},{9'b101110010},{9'b000100110},{9'b011001011},{9'b001010100},{9'b000100011},{9'b110011011},{9'b101111010},{9'b110101010},{9'b101001100},{9'b011101101},{9'b000001010},{9'b011000111},{9'b101111100},{9'b010101101},{9'b011110010},{9'b011000110},{9'b111101000},{9'b111111111},{9'b101110110},{9'b111010001},{9'b011000110},{9'b110100110},{9'b111011111},{9'b101000001},{9'b011111110},{9'b010110100},{9'b110100001},{9'b010001111},{9'b011011011},{9'b100010111},{9'b010110111},{9'b100001110},{9'b110100010},{9'b011001111},{9'b000100000},{9'b111000110},{9'b010100111},{9'b010111001},{9'b110100001},{9'b111001101},{9'b011100111},{9'b100010001},{9'b110101011},{9'b011011001},{9'b101001000},{9'b011000001},{9'b100000010},{9'b101110110},{9'b111111011},{9'b111000011},{9'b101010000},{9'b100100001},{9'b100110111},{9'b000100010},{9'b010000100},{9'b001101100},{9'b110011111},{9'b001000111},{9'b001101000},{9'b000001111},{9'b111111110},{9'b111101001},{9'b011111100},{9'b110010000},{9'b110010110},{9'b100000000},{9'b011000001},{9'b111000011},{9'b010110001},{9'b100000111},{9'b011010011},{9'b011011110},{9'b011001111},{9'b001010000},{9'b011100100},{9'b110011010},{9'b001101000},{9'b100010101},{9'b110011010},{9'b000101011},{9'b100110011},{9'b011100010},{9'b111001000},{9'b010000011},{9'b110011111},{9'b111101101},{9'b011101110},{9'b111000001},{9'b110111001},{9'b001111011},{9'b100000101},{9'b110011100},{9'b000011011},{9'b011001111},{9'b001000000},{9'b111111000},{9'b101111010},{9'b110000000},{9'b101101111},{9'b000010111},{9'b101011000},{9'b101011010},{9'b101011011},{9'b111011110},{9'b111100110},{9'b110000010},{9'b110100001},{9'b111000100},{9'b000000100},{9'b111010101},{9'b101000110},{9'b100010110},{9'b000110001},{9'b000011111},{9'b001001010},{9'b001011001},{9'b011100000},{9'b010000000},{9'b100111001},{9'b010010110},{9'b001110110},{9'b011010110},{9'b110010111},{9'b010001111},{9'b111101011},{9'b111111000},{9'b100111110},{9'b001100011},{9'b110111100},{9'b011110110},{9'b010010000},{9'b011011001},{9'b010011110},{9'b000111011},{9'b000101000},{9'b100110101},{9'b000101100},{9'b110011100},{9'b001101110},{9'b011010011},{9'b001111010},{9'b100111100},{9'b010110010},{9'b111011010},{9'b010011110},{9'b000111100},{9'b000100011},{9'b000011110},{9'b010011010},{9'b000111011},{9'b001001001},{9'b001011100},{9'b000011001},{9'b001000100},{9'b100000000},{9'b111101001},{9'b111000111},{9'b101000111},{9'b100110000},{9'b001100101},{9'b110001101},{9'b110010110},{9'b101001010},{9'b101001101},{9'b101001001},{9'b000010000},{9'b110101001},{9'b111000101},{9'b011101011},{9'b110100011},{9'b010011101},{9'b101010000},{9'b001001101},{9'b010111000},{9'b011110110},{9'b000101111},{9'b111110001},{9'b001010001},{9'b001001110},{9'b010011010},{9'b101101110},{9'b101111001},{9'b000011110},{9'b111111001},{9'b100001001},{9'b100101011},{9'b001001100},{9'b110001111},{9'b010111001},{9'b111100010},{9'b000111101},{9'b111100111},{9'b100111100},{9'b110010100},{9'b011000110},{9'b111000010},{9'b001110100},{9'b100111100},{9'b010100110},{9'b010011011},{9'b111011011},{9'b100110010},{9'b000010100},{9'b101010000},{9'b000010010},{9'b110001101},{9'b010011110},{9'b110010110},{9'b110110010},{9'b000110111},{9'b101101101},{9'b011010001},{9'b111001101},{9'b110000111},{9'b111100111},{9'b100001101},{9'b000111101},{9'b000101100},{9'b110100110},{9'b001110101},{9'b010000111},{9'b111000101},{9'b111101011},{9'b101000101},{9'b110011001},{9'b111101111},{9'b111100101},{9'b101011110},{9'b011010000},{9'b010111001},{9'b100010011},{9'b010110100},{9'b001100101},{9'b011010000},{9'b011011011},{9'b110011101},{9'b101100011},{9'b001010111},{9'b010100000},{9'b000101011},{9'b010111110},{9'b010011000},{9'b100110110},{9'b001000010},{9'b110000110},{9'b110001010},{9'b010000010},{9'b000001100},{9'b100011111},{9'b011110100},{9'b111011101},{9'b010010011},{9'b111111100},{9'b101101100},{9'b111010001},{9'b010010110},{9'b010011001},{9'b100101101},{9'b100001011},{9'b000111110},{9'b010010100},{9'b101111110},{9'b011001011},{9'b011001101},{9'b110000100},{9'b101001100},{9'b000000000},{9'b101101111},{9'b000001100},{9'b100011000},{9'b100011001},{9'b100001100},{9'b100000011},{9'b000100011},{9'b011100001},{9'b010101100},{9'b110111111},{9'b001010011},{9'b010100011},{9'b100111001},{9'b000110101},{9'b111010110},{9'b110111110},{9'b110001001},{9'b011101101},{9'b101010010},{9'b011011011},{9'b000101011},{9'b111000100},{9'b011001000},{9'b010100100},{9'b011110110},{9'b110111111},{9'b010010011},{9'b100000001},{9'b111000100},{9'b011100111},{9'b111111000},{9'b110001111},{9'b011010011},{9'b001011100},{9'b110010001},{9'b111001110},{9'b101110001},{9'b110001000},{9'b111000100},{9'b110001000},{9'b010101001},{9'b000111110},{9'b101111011},{9'b100001111},{9'b001111001},{9'b100010011},{9'b001000011},{9'b100101100},{9'b100010010},{9'b110010001},{9'b110001010},{9'b101000010},{9'b101101100},{9'b011110011},{9'b111000100},{9'b101001101},{9'b010111010},{9'b111000011},{9'b011101100},{9'b101001111},{9'b101001001},{9'b110100111},{9'b111111001},{9'b010100111},{9'b010111000},{9'b100001010},{9'b111111101},{9'b100001011},{9'b111100111},{9'b010001110},{9'b011001000},{9'b111111001},{9'b100000011},{9'b011001100},{9'b010100111},{9'b010011101},{9'b101100110},{9'b000000111},{9'b010110000},{9'b110111110},{9'b001000101},{9'b011101101},{9'b101100110},{9'b101100000},{9'b101110100},{9'b110001011},{9'b100011101},{9'b101101111},{9'b000011001},{9'b101000100},{9'b101111011},{9'b100100000},{9'b110111100},{9'b001110101},{9'b110010000},{9'b110001001},{9'b001111100},{9'b101010011},{9'b110000110},{9'b101110101},{9'b110001010},{9'b000001100},{9'b111111100},{9'b110111111},{9'b011110110},{9'b001111110},{9'b011111011},{9'b011011111},{9'b110110001},{9'b101000011},{9'b100110011},{9'b000110100},{9'b000011101},{9'b110000000},{9'b100110011},{9'b100010110},{9'b101110010},{9'b010011100},{9'b110011110},{9'b000101111},{9'b000001001},{9'b110100110},{9'b001010111},{9'b001011100},{9'b111100001},{9'b010101111},{9'b111110010},{9'b011111110},{9'b111101101},{9'b100000000},{9'b110011110},{9'b100011010},{9'b111111001},{9'b111000111},{9'b100000101},{9'b000110011},{9'b111101111},{9'b000010100},{9'b101101010},{9'b100100011},{9'b010011001},{9'b111110011},{9'b010000010},{9'b111010001},{9'b100110110},{9'b000111010},{9'b110111011},{9'b011100110},{9'b000001101},{9'b101100010},{9'b001100101},{9'b011010100},{9'b111100110},{9'b010011000},{9'b010000111},{9'b001011101},{9'b000000001},{9'b000010101},{9'b001111110},{9'b100111101},{9'b001101010},{9'b010110011},{9'b111000111},{9'b011111100},{9'b110011011},{9'b001100101},{9'b001010000},{9'b100110110},{9'b001111000},{9'b000100110},{9'b000101011},{9'b100011000},{9'b000110001},{9'b100000011},{9'b101010001},{9'b100101100},{9'b100000000},{9'b110110111},{9'b101001010},{9'b001110000},{9'b011000101},{9'b011101101},{9'b110110110},{9'b000001101},{9'b110011011},{9'b101100000},{9'b000111101},{9'b010100100},{9'b111111100},{9'b001001010},{9'b110101001},{9'b100101000},{9'b100011101},{9'b010100000},{9'b110101101},{9'b101101100},{9'b101011011},{9'b010000110},{9'b100000111},{9'b110100001},{9'b100111110},{9'b000001010},{9'b001011001},{9'b001100011},{9'b011110001},{9'b111100111},{9'b111111110},{9'b100000001},{9'b100011010},{9'b001111010},{9'b011111010},{9'b010000000},{9'b110111000},{9'b101011110},{9'b100010010},{9'b110011100},{9'b010011001},{9'b100101100},{9'b001101001},{9'b110000011},{9'b110011110},{9'b011100001},{9'b100010000},{9'b011001010},{9'b101010011},{9'b000010100},{9'b111010000},{9'b111110111},{9'b001110011},{9'b111001001},{9'b110110101},{9'b111101001},{9'b110100000},{9'b001010000},{9'b000110001},{9'b000111001},{9'b000001100},{9'b110110001},{9'b101100100},{9'b110110100},{9'b011001000},{9'b100010111},{9'b001001111},{9'b000100111},{9'b000111111},{9'b011011001},{9'b100011100},{9'b101001111},{9'b101111100},{9'b111001000},{9'b101000011},{9'b010000111},{9'b010001011},{9'b010010011},{9'b001000011},{9'b111000010},{9'b010011000},{9'b100010111},{9'b111101101},{9'b101100101},{9'b011001101},{9'b100100111},{9'b001110000},{9'b011001100},{9'b000001100},{9'b110011100},{9'b011001101},{9'b110010110},{9'b011011100},{9'b100110001},{9'b011100110},{9'b011100000},{9'b010110011},{9'b011100100},{9'b110110010},{9'b110001000},{9'b111011000},{9'b100011111},{9'b011000011},{9'b111001110},{9'b000011000},{9'b100101100},{9'b101100100},{9'b011001100},{9'b011101101},{9'b001010001},{9'b101000010},{9'b101101011},{9'b101001100},{9'b011011000},{9'b001110100},{9'b001101111},{9'b001100000},{9'b011100001},{9'b100000100},{9'b111001001},{9'b101000000},{9'b000110011},{9'b010101011},{9'b111010011},{9'b001110001},{9'b110000111},{9'b001110100},{9'b100101101},{9'b111110000},{9'b101000111},{9'b001100111},{9'b100011011},{9'b000111101},{9'b010001001},{9'b011001110},{9'b010001101},{9'b110101000},{9'b010110101},{9'b000101100},{9'b011100000},{9'b011011001},{9'b001001011},{9'b001000111},{9'b000100100},{9'b101100010},{9'b000011000},{9'b101011110},{9'b010011011},{9'b110110100},{9'b110001110},{9'b000110110},{9'b001110011},{9'b100111100},{9'b010011011},{9'b101001111},{9'b011001000},{9'b001000111},{9'b010100001},{9'b000010001},{9'b100100111},{9'b101000101},{9'b000010011},{9'b000001101},{9'b001001111},{9'b110001100},{9'b100000011},{9'b000000000},{9'b001110101},{9'b110101010},{9'b111010100},{9'b111010010},{9'b000111000},{9'b101101111},{9'b001101111},{9'b011110110},{9'b001110100},{9'b110010100},{9'b100111010},{9'b011010000},{9'b000001011},{9'b101100000},{9'b110011001},{9'b100001000},{9'b111001001},{9'b111000110},{9'b001111110},{9'b111101011},{9'b101011111},{9'b111110100},{9'b100101000},{9'b100100101},{9'b011000110},{9'b000010111},{9'b010111111},{9'b110101111},{9'b110111000},{9'b010010100},{9'b010010010},{9'b100100000},{9'b000001101},{9'b110001010},{9'b000110101},{9'b100101110},{9'b111100000},{9'b110011010},{9'b110001011},{9'b001000110},{9'b111000101},{9'b100111001},{9'b100010111},{9'b101100000},{9'b101001101},{9'b011000101},{9'b100001111},{9'b011101010},{9'b110111010},{9'b100001100},{9'b010011110},{9'b001101011},{9'b011011011},{9'b110000000},{9'b011110001},{9'b011101110},{9'b001000101},{9'b011111100},{9'b111100011},{9'b101110111},{9'b010001100},{9'b110001000},{9'b100111101},{9'b001001001},{9'b001100110},{9'b000110111},{9'b110110100},{9'b101010000},{9'b110100000},{9'b111010100},{9'b001100111},{9'b100010001},{9'b010001001},{9'b000111001},{9'b001000100},{9'b111001100},{9'b101010111},{9'b011110111},{9'b000100110},{9'b001100001},{9'b011101001},{9'b110110001},{9'b001001001},{9'b101110001},{9'b010011001},{9'b111011110},{9'b110111110},{9'b010011110},{9'b000100100},{9'b100011001},{9'b101010101},{9'b001101000},{9'b001100010},{9'b011001011},{9'b101101110},{9'b010110111},{9'b100111111},{9'b001101010},{9'b100111110},{9'b111000001},{9'b011101000},{9'b011001101},{9'b011000010},{9'b110101111},{9'b100011111},{9'b011001010},{9'b111110111},{9'b001100111},{9'b100100100},{9'b101001000},{9'b010110010},{9'b101000000},{9'b000010010},{9'b000001111},{9'b110101101},{9'b000101100},{9'b110011000},{9'b000000000},{9'b111011001},{9'b011110000},{9'b101100110},{9'b011000101},{9'b110100101},{9'b101010000},{9'b000100000},{9'b111011000},{9'b101111011},{9'b010111000},{9'b000100100},{9'b110100110},{9'b100101011},{9'b001111000},{9'b110110001},{9'b111111000},{9'b001100100},{9'b100011010},{9'b010011010},{9'b001010011},{9'b101001000},{9'b111110010},{9'b110000011},{9'b001100010},{9'b111011001},{9'b111000110},{9'b101001000},{9'b101001000},{9'b001101000},{9'b100110011},{9'b100011000},{9'b001000100},{9'b110010000},{9'b011110110},{9'b110100100},{9'b100010110},{9'b000111111},{9'b101000111},{9'b101110110},{9'b100100101},{9'b111001001},{9'b100011011},{9'b001100111},{9'b000001011},{9'b100111011},{9'b110001001},{9'b100111111},{9'b000001100},{9'b110110111},{9'b110110101},{9'b100000101},{9'b010100011},{9'b011101100},{9'b000100111},{9'b110100110},{9'b101011010},{9'b100111011},{9'b011100010},{9'b111001100},{9'b010001011},{9'b001010100},{9'b110001001},{9'b101110010},{9'b101010011},{9'b101110101},{9'b000110000},{9'b110010010},{9'b100001100},{9'b001111010},{9'b100011001},{9'b010000011},{9'b100010111},{9'b110111110},{9'b011001011},{9'b000100110},{9'b010000001},{9'b110100111},{9'b100000000},{9'b111010111},{9'b000110101},{9'b100100001},{9'b011110101},{9'b110011110},{9'b111101010},{9'b010101000},{9'b111000011},{9'b111100110},{9'b100110010},{9'b011000000},{9'b101000101},{9'b100100111},{9'b100101011},{9'b111100001},{9'b000001110},{9'b011000101},{9'b100100010},{9'b101101111},{9'b110011011},{9'b110111011},{9'b011101111},{9'b001111101},{9'b100111011},{9'b111000100},{9'b010011100},{9'b110000010},{9'b100101101},{9'b000010110},{9'b000010000},{9'b000001000},{9'b100001011},{9'b110111110},{9'b011011001},{9'b000110101},{9'b001001100},{9'b101000101},{9'b110111011},{9'b111001100},{9'b000100111},{9'b110100110},{9'b011100011},{9'b100000011},{9'b111100010},{9'b111111001},{9'b000100111},{9'b010111000},{9'b001011101},{9'b001100010},{9'b111100110},{9'b010001110},{9'b001011001},{9'b011111001},{9'b000000011},{9'b010101101},{9'b100000100},{9'b101110111},{9'b001111001},{9'b101010001},{9'b001101001},{9'b101111001},{9'b101011110},{9'b100101001},{9'b011101101},{9'b111010000},{9'b010111101},{9'b001000111},{9'b000010000},{9'b001010010},{9'b011011001},{9'b100100000},{9'b010001110},{9'b011110001},{9'b111111100},{9'b101000110},{9'b101101000},{9'b001001001},{9'b101000011},{9'b011010000},{9'b010010010},{9'b101101010},{9'b011101010},{9'b111101100},{9'b011111010},{9'b010011010},{9'b010001100},{9'b100110010},{9'b100000000},{9'b000101101},{9'b100101100},{9'b001000010},{9'b100001011},{9'b011100010},{9'b010010100},{9'b001101000},{9'b110001010},{9'b110010111},{9'b010111101},{9'b000101100},{9'b100011100},{9'b001110010},{9'b000011111},{9'b011111100},{9'b000100101},{9'b001000100},{9'b100011001},{9'b000001011},{9'b101010110},{9'b101000010},{9'b010011010},{9'b001111100},{9'b001110100},{9'b101110011},{9'b000110010},{9'b110010011},{9'b100110000},{9'b011000011},{9'b010100010},{9'b010111100},{9'b100110000},{9'b100000010},{9'b011111100},{9'b000100111},{9'b110111000},{9'b011011001},{9'b010101000},{9'b100101010},{9'b111011000},{9'b001100001},{9'b101010001},{9'b010011101},{9'b111011011},{9'b110101111},{9'b000100110},{9'b001001011},{9'b110100000},{9'b000111000},{9'b010011111},{9'b100110100},{9'b010011111},{9'b101011100},{9'b010011111},{9'b101011100},{9'b111000111},{9'b010100100},{9'b100101110},{9'b101101000},{9'b110011011},{9'b001011111},{9'b001101100},{9'b011101000},{9'b001111110},{9'b111011101},{9'b010110000},{9'b110101001},{9'b010011010},{9'b011100000},{9'b110001011},{9'b101000000},{9'b000001001},{9'b111100100},{9'b001101101},{9'b110111110},{9'b010111111},{9'b010111011},{9'b101000111},{9'b011111111},{9'b010101100},{9'b011010010},{9'b001101000},{9'b000011110},{9'b011001110},{9'b100101011},{9'b110011111},{9'b011010010},{9'b010111100},{9'b100110101},{9'b000001110},{9'b001110100},{9'b001101111},{9'b111101110},{9'b000111001},{9'b011110001},{9'b100001101},{9'b011001000},{9'b100011100},{9'b101110100},{9'b001000000},{9'b100011010},{9'b011000101},{9'b110111010},{9'b110101101},{9'b100100010},{9'b111000100},{9'b010100101},{9'b111101001},{9'b110011111},{9'b001011010},{9'b011010001},{9'b110010101},{9'b100100011},{9'b111001110},{9'b010101110},{9'b010011001},{9'b111110100},{9'b110101011},{9'b000111000},{9'b001110111},{9'b000001100},{9'b101101000},{9'b101001011},{9'b010011011},{9'b000000011},{9'b110100000},{9'b100001110},{9'b001110111},{9'b101001111},{9'b000111111},{9'b101010010},{9'b011110010},{9'b011000001},{9'b111011011},{9'b101100000},{9'b100000000},{9'b110100101},{9'b000011001},{9'b110101100},{9'b111010010},{9'b010100011},{9'b100101101},{9'b111011111},{9'b010111111},{9'b001110110},{9'b010110110},{9'b010111101},{9'b000101000},{9'b000001001},{9'b111001100},{9'b001000110},{9'b010000010},{9'b111001011},{9'b100110011},{9'b110000010},{9'b101110000},{9'b110001001},{9'b011101010},{9'b010111100},{9'b110110000},{9'b101011001},{9'b111000001},{9'b111011000},{9'b001101100},{9'b001110101},{9'b000011111},{9'b010011000},{9'b010110111},{9'b011000100},{9'b010111000},{9'b101110011},{9'b100001001},{9'b011111101},{9'b000111011},{9'b110100100},{9'b111000000},{9'b110100010},{9'b011101101},{9'b111101101},{9'b011010101},{9'b100100001},{9'b001101011},{9'b001111000},{9'b101010001},{9'b010111101},{9'b111101010},{9'b111100011},{9'b100010011},{9'b000110101},{9'b000101100},{9'b011101011},{9'b100010010},{9'b110011101},{9'b010100101},{9'b111000001},{9'b100001000},{9'b100011010},{9'b001000001},{9'b110101011},{9'b011001010},{9'b111010010},{9'b111100000},{9'b000001100},{9'b010111011},{9'b010001111},{9'b010101111},{9'b110000110},{9'b011110111},{9'b111011100},{9'b101100110},{9'b010000001},{9'b010001110},{9'b101111100},{9'b000001010},{9'b010011011},{9'b011101101},{9'b011001010},{9'b011111100},{9'b011010101},{9'b011001111},{9'b001110111},{9'b100100001},{9'b101111000},{9'b111101011},{9'b010111010},{9'b110001000},{9'b011100010},{9'b101100101},{9'b100010001},{9'b101001100},{9'b110110000},{9'b110001011},{9'b101110100},{9'b000011000},{9'b100100011},{9'b100001001},{9'b110101100},{9'b001010001},{9'b100100110},{9'b110110000},{9'b010110100},{9'b000011011},{9'b111011101},{9'b111010111},{9'b100110110},{9'b001001100},{9'b010010011},{9'b110000100},{9'b010000110},{9'b010010010},{9'b000111100},{9'b000000100},{9'b011111111},{9'b011011101},{9'b010100101},{9'b000000010},{9'b111001111},{9'b110110111},{9'b111101011},{9'b000010100},{9'b011111000},{9'b010000110},{9'b000110101},{9'b111100100},{9'b101101011},{9'b001001100},{9'b001111001},{9'b110001011},{9'b110111101},{9'b111000100},{9'b111100101},{9'b110001111},{9'b010111100},{9'b111000011},{9'b011010101},{9'b100001001},{9'b100101111},{9'b100111111},{9'b111010110},{9'b101101000},{9'b000000100},{9'b001000101},{9'b010010010},{9'b000001111},{9'b011100001},{9'b000100001},{9'b001010100},{9'b000001000},{9'b000010111},{9'b110001111},{9'b111000010},{9'b011001011},{9'b111110101},{9'b100001100},{9'b010011010},{9'b010110100},{9'b011110100},{9'b010111100},{9'b000010100},{9'b000111111},{9'b101101011},{9'b101011100},{9'b011011111},{9'b000111101},{9'b010001000},{9'b100010101},{9'b000111110},{9'b010110001},{9'b111001010},{9'b100111001},{9'b001111000},{9'b001110111},{9'b000001001},{9'b100101110},{9'b111111011},{9'b110010011},{9'b110000111},{9'b111101110},{9'b001101110},{9'b001111110},{9'b110111101},{9'b000110101},{9'b101111101},{9'b010001100},{9'b100001110},{9'b101111001},{9'b111101000},{9'b001001010},{9'b011110000},{9'b101110110},{9'b110001101},{9'b100010000},{9'b111110101},{9'b110110000},{9'b010000000},{9'b111000010},{9'b000111101},{9'b100011111},{9'b111000011},{9'b100010110},{9'b111101000},{9'b000100011},{9'b110011101},{9'b100011110},{9'b001100001},{9'b100001100},{9'b110000000},{9'b001101011},{9'b011100110},{9'b000101000},{9'b011010100},{9'b100000011},{9'b000101000},{9'b000101100},{9'b011000010},{9'b000010001},{9'b011010011},{9'b010011100},{9'b100100111},{9'b100001001},{9'b101010001},{9'b100011100},{9'b011000111},{9'b110101010},{9'b110111001},{9'b101000101},{9'b101100011},{9'b101000100},{9'b011010101},{9'b001011001},{9'b011000101},{9'b100100011},{9'b101011111},{9'b001000010},{9'b111010101},{9'b011000011},{9'b001111001},{9'b111101000},{9'b011011001},{9'b010001011},{9'b101010010},{9'b000110010},{9'b101110011},{9'b111000000},{9'b001010010},{9'b101001000},{9'b010111010},{9'b101100011},{9'b111011110},{9'b000010111},{9'b111001010},{9'b011000111},{9'b101110010},{9'b101100100},{9'b110000100},{9'b000010101},{9'b011110111},{9'b010000111},{9'b110111110},{9'b100010100},{9'b011001001},{9'b001111101},{9'b001100101},{9'b100001111},{9'b101111000},{9'b110010010},{9'b110101100},{9'b100011001},{9'b101100101},{9'b001000000},{9'b110111010},{9'b000001101},{9'b011110001},{9'b110110101},{9'b010010001},{9'b001000101},{9'b111011001},{9'b111000101},{9'b111111000},{9'b010001101},{9'b011110111},{9'b000000110},{9'b011011000},{9'b010000000},{9'b001110010},{9'b110111000},{9'b000010100},{9'b011100101},{9'b101101110},{9'b110101100},{9'b011100011},{9'b111001000},{9'b001110110},{9'b110010111},{9'b110111111},{9'b001110101},{9'b101100011},{9'b110101101},{9'b101111111},{9'b001011010},{9'b101100101},{9'b110011011},{9'b010111001},{9'b000001111},{9'b011111001},{9'b011101000},{9'b001101000},{9'b110011100},{9'b111001100},{9'b000111100},{9'b100100101},{9'b011000101},{9'b011001101},{9'b110001010},{9'b111001000},{9'b101100110},{9'b011001001},{9'b001000000},{9'b010011011},{9'b010111000},{9'b100110001},{9'b100100101},{9'b111110000},{9'b111001111},{9'b100011011},{9'b110011010},{9'b111111111},{9'b101101000},{9'b100000010},{9'b110100001},{9'b011000111},{9'b111100010},{9'b111000011},{9'b001000010},{9'b010101011},{9'b110010010},{9'b010101011},{9'b110111100},{9'b100001111},{9'b010111001},{9'b110010001},{9'b101100011},{9'b011111001},{9'b011001010},{9'b100000000},{9'b101010111},{9'b010011000},{9'b000101110},{9'b001110100},{9'b010100110},{9'b010011011},{9'b001101100},{9'b010010001},{9'b010110100},{9'b010111000},{9'b111100011},{9'b011000011},{9'b001100110},{9'b101011101},{9'b011000001},{9'b101000010},{9'b101110011},{9'b010000001},{9'b110000001},{9'b010011011},{9'b111001110},{9'b111101110},{9'b011110000},{9'b011010101},{9'b001100100},{9'b001100011},{9'b111011100},{9'b100000110},{9'b010110011},{9'b011101111},{9'b111001001},{9'b100111110},{9'b001110000},{9'b010101111},{9'b011001001},{9'b100111010},{9'b111110000},{9'b000100100},{9'b001010000},{9'b101000101},{9'b010000000},{9'b011100000},{9'b111011001},{9'b100100110},{9'b111010111},{9'b010000110},{9'b101010000},{9'b011001011},{9'b100100110},{9'b000011010},{9'b001100000},{9'b100010001},{9'b001111101},{9'b010111011},{9'b110001011},{9'b001001001},{9'b110110111},{9'b011010001},{9'b010101011},{9'b110111111},{9'b101011010},{9'b111010011},{9'b100101000},{9'b010110101},{9'b110101000},{9'b111101101},{9'b110100100},{9'b010011000},{9'b010111000},{9'b001001111},{9'b000010100},{9'b101110011},{9'b010011101},{9'b110110011},{9'b101110011},{9'b110000000},{9'b101011000},{9'b101110001},{9'b111110010},{9'b000110110},{9'b000101101},{9'b110111111},{9'b010111101},{9'b011010101},{9'b010111100},{9'b110001000},{9'b000010101},{9'b101101101},{9'b100110100},{9'b001111010},{9'b111011110},{9'b100111110},{9'b011110001},{9'b011001001},{9'b110001101},{9'b111111110},{9'b010101000},{9'b000001011},{9'b001100100},{9'b101011111},{9'b011101110},{9'b110100111},{9'b111100000},{9'b110100101},{9'b110101000},{9'b010110001},{9'b111011011},{9'b100001001},{9'b111011101},{9'b100111101},{9'b001111110},{9'b000011010},{9'b111110011},{9'b101000000},{9'b000110010},{9'b111010011},{9'b100101111},{9'b100001110},{9'b100011011},{9'b110100010},{9'b000000111},{9'b011100111},{9'b000000110},{9'b101010001},{9'b100000011},{9'b000111001},{9'b011001000},{9'b001101111},{9'b100010111},{9'b000001110},{9'b110101100},{9'b110000011},{9'b111000111},{9'b011100111},{9'b110000101},{9'b100101011},{9'b001000101},{9'b001001101},{9'b110001010},{9'b010000000},{9'b111011010},{9'b110101110},{9'b011111000},{9'b101101000},{9'b010100110},{9'b011101010},{9'b111001101},{9'b010111011},{9'b001111100},{9'b110100011},{9'b001001000},{9'b100010101},{9'b001110100},{9'b001101001},{9'b001111100},{9'b110110101},{9'b011110001},{9'b100000000},{9'b001001010},{9'b110010010},{9'b001010101},{9'b111001110},{9'b011011011},{9'b001110000},{9'b100110000},{9'b010100100},{9'b001000011},{9'b000000000},{9'b110000010},{9'b001000001},{9'b001100000},{9'b011011000},{9'b001100100},{9'b011011011},{9'b100110111},{9'b000011010},{9'b011101011},{9'b101110100},{9'b100111011},{9'b001111011},{9'b111111000},{9'b101110110},{9'b111101011},{9'b001100001},{9'b010110010},{9'b110000111},{9'b010101000},{9'b010100010},{9'b011111010},{9'b001101110},{9'b011111010},{9'b100100010},{9'b100001101},{9'b001100101},{9'b000000011},{9'b101001011},{9'b100110100},{9'b101001111},{9'b001111000},{9'b011111101},{9'b101010000},{9'b111101010},{9'b101110110},{9'b101000111},{9'b100110010},{9'b000100001},{9'b111011111},{9'b111011010},{9'b000000010},{9'b001101000},{9'b111010101},{9'b100111001},{9'b111100000},{9'b011100010},{9'b111000000},{9'b010010110},{9'b100001011},{9'b100010101},{9'b111001001},{9'b001011010},{9'b101000010},{9'b010100000},{9'b100000110},{9'b101110000},{9'b001110100},{9'b011011011},{9'b111111100},{9'b111010010},{9'b100100100},{9'b110100110},{9'b111110111},{9'b011110001},{9'b001010101},{9'b111010010},{9'b111010110},{9'b111100011},{9'b010100011},{9'b010110001},{9'b010101000},{9'b011001000},{9'b011101000},{9'b111110100},{9'b111000111},{9'b110101101},{9'b110100001},{9'b010001111},{9'b001110101},{9'b110010011},{9'b111001110},{9'b000111100},{9'b000010000},{9'b101111001},{9'b111010100},{9'b000110011},{9'b101101000},{9'b100110110},{9'b110001000},{9'b001000011},{9'b001010001},{9'b110101001},{9'b010110101},{9'b101001101},{9'b101101110},{9'b001000010},{9'b100010100},{9'b110100011},{9'b001001110},{9'b001101111},{9'b100010100},{9'b110011010},{9'b110000100},{9'b100100110},{9'b111011001},{9'b000010001},{9'b010100001},{9'b010100011},{9'b000011101},{9'b101000100},{9'b101110100},{9'b010101101},{9'b101011000},{9'b100100011},{9'b000001100},{9'b011110011},{9'b011110101},{9'b011000011},{9'b011000010},{9'b110110010},{9'b001110001},{9'b011111110},{9'b000010001},{9'b000111001},{9'b110110011},{9'b001100100},{9'b000000011},{9'b111001111},{9'b111001110},{9'b100100111},{9'b011100000},{9'b101010010},{9'b101100101},{9'b111001001},{9'b011010110},{9'b010110101},{9'b001000111},{9'b010101000},{9'b011011011},{9'b010001101},{9'b010110010},{9'b001100001},{9'b001111000},{9'b000101000},{9'b011010111},{9'b101001010},{9'b101110100},{9'b100011111},{9'b011101110},{9'b010010101},{9'b001101001},{9'b110010010},{9'b101001010},{9'b010010010},{9'b110110011},{9'b111110100},{9'b010001000},{9'b010110101},{9'b001010011},{9'b101000110},{9'b110110101},{9'b011100110},{9'b110010101},{9'b100001011},{9'b011110000},{9'b010011101},{9'b001001111},{9'b010111001},{9'b100101101},{9'b110111111},{9'b101111011},{9'b111110000},{9'b011111001},{9'b001010001},{9'b001101001},{9'b100101111},{9'b000110110},{9'b001111111},{9'b000111100},{9'b100010010},{9'b000010101},{9'b011000011},{9'b011000011},{9'b101100010},{9'b010001110},{9'b101010001},{9'b010100001},{9'b000111110},{9'b001001001},{9'b101101101},{9'b000000101},{9'b000101110},{9'b111000011},{9'b001111101},{9'b101111000},{9'b010110000},{9'b011000110},{9'b010000110},{9'b101111110},{9'b101101110},{9'b111110111},{9'b100111010},{9'b010111000},{9'b000110110},{9'b111010111},{9'b100000111},{9'b111110000},{9'b110001001},{9'b001101100},{9'b100101111},{9'b110111001},{9'b010010101},{9'b001011110},{9'b101101100},{9'b101010110},{9'b010001001},{9'b110101111},{9'b001110010},{9'b011100000},{9'b010100010},{9'b111011100},{9'b001000010},{9'b110110111},{9'b100001011},{9'b100100110},{9'b011110000},{9'b000011111},{9'b011101100},{9'b000000011},{9'b001010111},{9'b010010001},{9'b110000010},{9'b001110010},{9'b111100100},{9'b110111100},{9'b000011011},{9'b101000110},{9'b100111110},{9'b111010110},{9'b101010110},{9'b111101010},{9'b110110100},{9'b001000011},{9'b010011101},{9'b110110100},{9'b111011101},{9'b100011100},{9'b100111001},{9'b000111111},{9'b110100110},{9'b011010100},{9'b101001010},{9'b111110100},{9'b111010100},{9'b000000111},{9'b111000110},{9'b100111100},{9'b010000001},{9'b101111011},{9'b011101111},{9'b011100101},{9'b000001011},{9'b011101010},{9'b111101001},{9'b010100011},{9'b011110000},{9'b001011001},{9'b000111011},{9'b011011101},{9'b101110001},{9'b000101111},{9'b001001100},{9'b101101111},{9'b010010001},{9'b100111101},{9'b111100101},{9'b011001001},{9'b100100100},{9'b001111100},{9'b111101011},{9'b111101011},{9'b001110010},{9'b000001000},{9'b011100001},{9'b010011111},{9'b111000100},{9'b010000110},{9'b100001011},{9'b101000111},{9'b001101100},{9'b000000000},{9'b001101000},{9'b011101111},{9'b010011110},{9'b011111011},{9'b111011011},{9'b100110100},{9'b000011011},{9'b000010000},{9'b111110010},{9'b011010111},{9'b001011111},{9'b001101100},{9'b100001101},{9'b101010000},{9'b011010010},{9'b101111000},{9'b100000010},{9'b011101010},{9'b100111011},{9'b011110010},{9'b110101100},{9'b100101000},{9'b101111100},{9'b000100101},{9'b011110100},{9'b111011011},{9'b001101111},{9'b001010111},{9'b011010000},{9'b010011111},{9'b000001000},{9'b101111000},{9'b111001101},{9'b100111100},{9'b001011101},{9'b001110011},{9'b110000000},{9'b111100100},{9'b111011110},{9'b101011111},{9'b001000111},{9'b110010001},{9'b110010010},{9'b000001111},{9'b010101010},{9'b010010110},{9'b101010011},{9'b011001101},{9'b001101101},{9'b011111001},{9'b011100100},{9'b001100100},{9'b111010001},{9'b101001010},{9'b011011000},{9'b101111111},{9'b011000100},{9'b110001001},{9'b110010010},{9'b011101010},{9'b100010100},{9'b011001100},{9'b011100101},{9'b110101011},{9'b101111000},{9'b000010011},{9'b010001100},{9'b001111101},{9'b100100000},{9'b110101011},{9'b010110010},{9'b011010001},{9'b111010010},{9'b111110001},{9'b110111010},{9'b011110101},{9'b110001100},{9'b000011011},{9'b000011111},{9'b101111011},{9'b100101011},{9'b110011001},{9'b110001011},{9'b110001110},{9'b110101010},{9'b100100000},{9'b001111100},{9'b100100101},{9'b010110100},{9'b110011001},{9'b011101011},{9'b101110010},{9'b001010110},{9'b010011110},{9'b010000011},{9'b011011101},{9'b101000111},{9'b101110111},{9'b100011101},{9'b110010000},{9'b100101100},{9'b011100010},{9'b111101101},{9'b101111001},{9'b000000111},{9'b010010101},{9'b100010010},{9'b100001100},{9'b101101001},{9'b100111010},{9'b110110100},{9'b100110001},{9'b111000010},{9'b101111010},{9'b101110110},{9'b110000000},{9'b010101100},{9'b100111100},{9'b111001110},{9'b101001001},{9'b010001001},{9'b010001010},{9'b111000101},{9'b100010111},{9'b101011100},{9'b111010011},{9'b111011000},{9'b000110111},{9'b110000101},{9'b111100000},{9'b111001010},{9'b110000100},{9'b011011001},{9'b101011011},{9'b111010011},{9'b000010000},{9'b000100110},{9'b100010010},{9'b111111101},{9'b000110010},{9'b011111110},{9'b100011101},{9'b100100001},{9'b010110001},{9'b000001100},{9'b111001000},{9'b100110110},{9'b010000010},{9'b010101110},{9'b101110001},{9'b001001111},{9'b000001001},{9'b011110000},{9'b110010110},{9'b011101001},{9'b101001101},{9'b100111000},{9'b101100110},{9'b001111101},{9'b101011010},{9'b010101001},{9'b001111100},{9'b001000011},{9'b010001000},{9'b010100111},{9'b001101001},{9'b110010001},{9'b010110010},{9'b100011000},{9'b110010011},{9'b101110111},{9'b101011010},{9'b001111011},{9'b100101001},{9'b000011100},{9'b100110000},{9'b111111001},{9'b110110011},{9'b100011100},{9'b000101100},{9'b110010101},{9'b001001001},{9'b011111100},{9'b111111001},{9'b001001101},{9'b000100010},{9'b100011001},{9'b100001110},{9'b110011010},{9'b111010110},{9'b001100011},{9'b101111110},{9'b001011001},{9'b111001110},{9'b000011011},{9'b001101000},{9'b000101010},{9'b101101001},{9'b110110001},{9'b000100010},{9'b010001010},{9'b000010110},{9'b111011101},{9'b000111011},{9'b110111000},{9'b000010101},{9'b001000010},{9'b111001100},{9'b001110010},{9'b111000011},{9'b001100000},{9'b011110001},{9'b000000100},{9'b100000110},{9'b000111100},{9'b110110111},{9'b010110101},{9'b110011011},{9'b001101011},{9'b111111100},{9'b110111111},{9'b001110010},{9'b101101100},{9'b100110010},{9'b010110010},{9'b101011100},{9'b101111111},{9'b000100011},{9'b001101100},{9'b110010001},{9'b101010000},{9'b100000011},{9'b001100011},{9'b111001101},{9'b111011100},{9'b000000111},{9'b000110101},{9'b011111110},{9'b001010011},{9'b010000111},{9'b011100000},{9'b001000001},{9'b010000100},{9'b100000001},{9'b101001011},{9'b100010001},{9'b001100010},{9'b000110100},{9'b011111100},{9'b010011011},{9'b110100000},{9'b001110101},{9'b100011100},{9'b100100111},{9'b010010000},{9'b001001110},{9'b001011100},{9'b010000010},{9'b010111011},{9'b100100101},{9'b010000011},{9'b001011000},{9'b001110101},{9'b100100000},{9'b011010010},{9'b111001101},{9'b111000100},{9'b001111100},{9'b110101111},{9'b010001010},{9'b000001000},{9'b001111001},{9'b101000111},{9'b111111110},{9'b100111110},{9'b011110110},{9'b110011110},{9'b001110000},{9'b011111110},{9'b000011000},{9'b010110000},{9'b100011000},{9'b011100001},{9'b011010111},{9'b011010000},{9'b010110111},{9'b000000010},{9'b101111000},{9'b101001101},{9'b100110100},{9'b010010001},{9'b011111111},{9'b111100100},{9'b011100010},{9'b111100000},{9'b100011001},{9'b000100010},{9'b101011110},{9'b010011100},{9'b010000100},{9'b001110100},{9'b101110001},{9'b101001011},{9'b101010111},{9'b110000101},{9'b011100110},{9'b100010100},{9'b000011011},{9'b000100011},{9'b111110101},{9'b110100111},{9'b110001111},{9'b110010001},{9'b111110101},{9'b000110110},{9'b011001010},{9'b010100111},{9'b001001100},{9'b011011010},{9'b110101010},{9'b001100001},{9'b100101100},{9'b011110100},{9'b111111110},{9'b111100110},{9'b100100011},{9'b000110011},{9'b010000111},{9'b111110010},{9'b010010101},{9'b111010111},{9'b001101100},{9'b110101110},{9'b100110110},{9'b000111100},{9'b100110110},{9'b010011101},{9'b110010100},{9'b111001111},{9'b100001011},{9'b100101100},{9'b010100001},{9'b111101110},{9'b010010001},{9'b001011000},{9'b101010101},{9'b011100100},{9'b000111010},{9'b100111011},{9'b001000001},{9'b111101111},{9'b110100111},{9'b010111010},{9'b011000011},{9'b110000100},{9'b100010100},{9'b110110001},{9'b000110110},{9'b110101100},{9'b001011100},{9'b100000100},{9'b011011010},{9'b111110011},{9'b001001011},{9'b011000001},{9'b111110110},{9'b101010111},{9'b011101001},{9'b000010111},{9'b010010110},{9'b111000101},{9'b000011001},{9'b001111011},{9'b111110101},{9'b110101010},{9'b011110001},{9'b010111111},{9'b010111011},{9'b110010100},{9'b011110111},{9'b101000111},{9'b011000110},{9'b010100000},{9'b000010101},{9'b111011111},{9'b111100010},{9'b111011010},{9'b100000101},{9'b110010001},{9'b010101100},{9'b101011110},{9'b101010110},{9'b000000111},{9'b100001110},{9'b011101111},{9'b110010001},{9'b010111010},{9'b011100011},{9'b101110110},{9'b101001001},{9'b111101010},{9'b110101100},{9'b010011010},{9'b101101101},{9'b011111110},{9'b010010001},{9'b001111011},{9'b110101010},{9'b111110100},{9'b110001001},{9'b110101101},{9'b111110011},{9'b000110100},{9'b010100101},{9'b001100101},{9'b110001111},{9'b011110010},{9'b011000010},{9'b100010010},{9'b010010000},{9'b010001001},{9'b101111100},{9'b110100101},{9'b011011111},{9'b110001100},{9'b011101100},{9'b110111001},{9'b011001011},{9'b011110000},{9'b010010001},{9'b111011000},{9'b001111110},{9'b101101101},{9'b111001001},{9'b011011001},{9'b111011010},{9'b101111011},{9'b000110000},{9'b100101111},{9'b000000000},{9'b110100101},{9'b101000001},{9'b011000101},{9'b111000010},{9'b110001101},{9'b100010011},{9'b010011100},{9'b001010111},{9'b101001111},{9'b111101011},{9'b000111010},{9'b010110010},{9'b001100001},{9'b101110000},{9'b100100100},{9'b100001101},{9'b010000011},{9'b100001101},{9'b111011000},{9'b111001100},{9'b011000111},{9'b010000100},{9'b011000011},{9'b101011000},{9'b110110110},{9'b101100101},{9'b001101100},{9'b000100110},{9'b001011010},{9'b011010011},{9'b000101101},{9'b011011010},{9'b001011110},{9'b000000000},{9'b110010011},{9'b110101001},{9'b110101111},{9'b101010110},{9'b111100011},{9'b100100001},{9'b110111111},{9'b011001011},{9'b111000101},{9'b110011111},{9'b111100010},{9'b010110010},{9'b110010110},{9'b101000000},{9'b101100101},{9'b000101111},{9'b000111101},{9'b111000110},{9'b000111010},{9'b101100001},{9'b101001011},{9'b101101100},{9'b111010101},{9'b101000011},{9'b010011100},{9'b110001110},{9'b101100011},{9'b001000010},{9'b001001000},{9'b001001001},{9'b001100001},{9'b101001010},{9'b010110100},{9'b010001011},{9'b110001101},{9'b101101000},{9'b010011011},{9'b011011010},{9'b010110101},{9'b111110110},{9'b111010101},{9'b111000110},{9'b001000011},{9'b100000110},{9'b110100011},{9'b110100100},{9'b111001001},{9'b000000110},{9'b100110100},{9'b100110111},{9'b110010101},{9'b100011110},{9'b000101111},{9'b100010100},{9'b000110111},{9'b110110101},{9'b011000101},{9'b100100001},{9'b001000011},{9'b010000010},{9'b000101000},{9'b110001111},{9'b010010100},{9'b001000000},{9'b010110011},{9'b010001001},{9'b000111111},{9'b111110011},{9'b001101011},{9'b100001001},{9'b010111011},{9'b011101001},{9'b100110010},{9'b010010100},{9'b111000001},{9'b010010100},{9'b111111101},{9'b111001001},{9'b101100111},{9'b000011100},{9'b001111001},{9'b111000010},{9'b001110110},{9'b100100001},{9'b101111001},{9'b001101101},{9'b001011101},{9'b111000001},{9'b010010000},{9'b111101101},{9'b101110101},{9'b000011110},{9'b000011100},{9'b100000111},{9'b100010110},{9'b111001000},{9'b000101010},{9'b110011011},{9'b111100011},{9'b101101101},{9'b110111101},{9'b011011111},{9'b111110110},{9'b110101011},{9'b010111000},{9'b011110010},{9'b111100000},{9'b001111110},{9'b010011110},{9'b111110111},{9'b000010001},{9'b101001100},{9'b101001110},{9'b111010101},{9'b001111011},{9'b101001010},{9'b000000011},{9'b000000001},{9'b001100101},{9'b000101111},{9'b010010011},{9'b111101100},{9'b110011110},{9'b000110101},{9'b110000010},{9'b000101001},{9'b001010010},{9'b110100100},{9'b110000001},{9'b110001011},{9'b100111011},{9'b111111110},{9'b101100111},{9'b101101001},{9'b010010011},{9'b011000011},{9'b111010100},{9'b101011101},{9'b111101011},{9'b000110000},{9'b110100110},{9'b101011100},{9'b101110001},{9'b110001001},{9'b010001011},{9'b111110101},{9'b101011000},{9'b011010010},{9'b110111110},{9'b110110010},{9'b000111010},{9'b101100011},{9'b011011100},{9'b111000110},{9'b101110001},{9'b100011100},{9'b000010111},{9'b010001001},{9'b011111101},{9'b000110010},{9'b110111000},{9'b000000110},{9'b111011110},{9'b000011111},{9'b010001001},{9'b000111011},{9'b000001000},{9'b000010000},{9'b111011110},{9'b010111011},{9'b001001010},{9'b011001111},{9'b101011100},{9'b000001110},{9'b001001101},{9'b000101000},{9'b101101011},{9'b100001010},{9'b001011001},{9'b010100100},{9'b010101111},{9'b000110011},{9'b011110110},{9'b001100101},{9'b000000011},{9'b100100010},{9'b110011011},{9'b011111100},{9'b111100011},{9'b001111110},{9'b001011010},{9'b100110110},{9'b111000110},{9'b000101100},{9'b111100100},{9'b100010010},{9'b011110001},{9'b100010011},{9'b110111100},{9'b100001100},{9'b101000100},{9'b110101111},{9'b111110011},{9'b001010101},{9'b110110110},{9'b100010001},{9'b111111111},{9'b011110011},{9'b101010000},{9'b010100011},{9'b110010100},{9'b011100010},{9'b111101000},{9'b001111111},{9'b101100110},{9'b001110101},{9'b111101010},{9'b000001001},{9'b011101000},{9'b111111101},{9'b100100101},{9'b101111000},{9'b001100011},{9'b111011110},{9'b011110010},{9'b110100000},{9'b100101001},{9'b101101100},{9'b000011100},{9'b001110000},{9'b010010111},{9'b111001101},{9'b001010011},{9'b110110100},{9'b000010010},{9'b001101110},{9'b100001001},{9'b111010001},{9'b110101011},{9'b000101000},{9'b011100001},{9'b001110010},{9'b110011111},{9'b010010101},{9'b010111111},{9'b100001000},{9'b110100110},{9'b010101101},{9'b011101011},{9'b000110011},{9'b001000011},{9'b111001011},{9'b000100100},{9'b111010111},{9'b110000111},{9'b101111101},{9'b000011001},{9'b110011011},{9'b000101110},{9'b111000001},{9'b101100101},{9'b101101011},{9'b001101011},{9'b111101111},{9'b110110101},{9'b110010101},{9'b111110100},{9'b010010010},{9'b110001110},{9'b101000001},{9'b101100000},{9'b111000101},{9'b010101101},{9'b000011111},{9'b011010001},{9'b100001111},{9'b000011010},{9'b000101101},{9'b000100110},{9'b001011000},{9'b101100000},{9'b000011011},{9'b010010000},{9'b111111110},{9'b000110110},{9'b100110010},{9'b010111011},{9'b110110101},{9'b001001100},{9'b101110111},{9'b001010011},{9'b100000010},{9'b110001110},{9'b010010001},{9'b101010111},{9'b000010100},{9'b111011100},{9'b011110101},{9'b000110110},{9'b100101001},{9'b011101000},{9'b101010101},{9'b000101001},{9'b101001111},{9'b001011111},{9'b100001011},{9'b101000110},{9'b010010111},{9'b010110111},{9'b001100010},{9'b110001110},{9'b001111010},{9'b011001001},{9'b110111101},{9'b110111110},{9'b000010100},{9'b001101010},{9'b000101100},{9'b101010000},{9'b110000000},{9'b111100001},{9'b100100100},{9'b011101100},{9'b100010110},{9'b111000011},{9'b101001110},{9'b101001110},{9'b000011001},{9'b000001100},{9'b010110010},{9'b010000100},{9'b001001000},{9'b011101001},{9'b011110011},{9'b010011001},{9'b010100111},{9'b011100111},{9'b110111000},{9'b100001011},{9'b100011001},{9'b010101110},{9'b110101010},{9'b101100111},{9'b101001001},{9'b010000111},{9'b111101010},{9'b110001001},{9'b000011000},{9'b100100110},{9'b110110010},{9'b010101110},{9'b111111011},{9'b111001110},{9'b101010100},{9'b011000110},{9'b101001011},{9'b111010001},{9'b000011011},{9'b011011001},{9'b101010111},{9'b011011110},{9'b110011001},{9'b010000100},{9'b110001010},{9'b111101010},{9'b110111011},{9'b110111000},{9'b101010001},{9'b000100001},{9'b111011010},{9'b110011100},{9'b011000111},{9'b111110110},{9'b001101001},{9'b100101110},{9'b110001011},{9'b000110000},{9'b010011111},{9'b011101100},{9'b111101011},{9'b110111100},{9'b110110111},{9'b001100101},{9'b011011001},{9'b010001110},{9'b000111111},{9'b000000000},{9'b100000001},{9'b010110100},{9'b010011110},{9'b011110000},{9'b011011010},{9'b111101011},{9'b010100010},{9'b001001011},{9'b101001010},{9'b000011100},{9'b001111110},{9'b111110000},{9'b011001111},{9'b000101001},{9'b000011110},{9'b000110100},{9'b111011100},{9'b101101000},{9'b101001111},{9'b100110101},{9'b100110110},{9'b100110110},{9'b001010010},{9'b001100100},{9'b010100110},{9'b001101011},{9'b000101010},{9'b011100010},{9'b010010100},{9'b000011110},{9'b110111011},{9'b111111010},{9'b001001000},{9'b101001101},{9'b011110110},{9'b110010100},{9'b001011010},{9'b001110110},{9'b011000111},{9'b100000111},{9'b000111110},{9'b010011101},{9'b010000111},{9'b111110110},{9'b010011100},{9'b001010101},{9'b100110110},{9'b110111010},{9'b011110001},{9'b110011110},{9'b001000001},{9'b111101110},{9'b101101011},{9'b011100010},{9'b011110111},{9'b001010010},{9'b111001100},{9'b010111100},{9'b011100111},{9'b011111001},{9'b100101101},{9'b000111001},{9'b001111001},{9'b010111011},{9'b111000010},{9'b100101110},{9'b110100111},{9'b010111011},{9'b001111010},{9'b110011010},{9'b111110010},{9'b000101110},{9'b011100111},{9'b110111000},{9'b110110011},{9'b010011111},{9'b111101011},{9'b110001110},{9'b011111011},{9'b011010001},{9'b101011111},{9'b001101010},{9'b110110100},{9'b110111011},{9'b010011000},{9'b111100100},{9'b010010011},{9'b111010001},{9'b010001101},{9'b101110000},{9'b111110010},{9'b010100010},{9'b101101101},{9'b100010110},{9'b011110111},{9'b110101001},{9'b001100101},{9'b101000110},{9'b010110000},{9'b110000001},{9'b001010011},{9'b001010100},{9'b111000110},{9'b100000110},{9'b000101010},{9'b111011001},{9'b001100000},{9'b000001100},{9'b101111110},{9'b110111001},{9'b100110010},{9'b010111001},{9'b101001011},{9'b001010011},{9'b110100000},{9'b001100100},{9'b010101010},{9'b011010011},{9'b011011100},{9'b101010010},{9'b001110101},{9'b111000110},{9'b001011001},{9'b101110000},{9'b101110010},{9'b110010000},{9'b101111110},{9'b001000100},{9'b001010010},{9'b011010001},{9'b100110110},{9'b100110100},{9'b101001001},{9'b110011100},{9'b111111111},{9'b111111111},{9'b100110101},{9'b110111100},{9'b110110101},{9'b011010111},{9'b100001111},{9'b001101011},{9'b101010000},{9'b100111110},{9'b001111110},{9'b111001101},{9'b101000111},{9'b000111111},{9'b010110000},{9'b101100100},{9'b101110011},{9'b101010000},{9'b111111110},{9'b000110101},{9'b000001110},{9'b101100011},{9'b111011101},{9'b010100110},{9'b110001010},{9'b110101011},{9'b101001000},{9'b011010011},{9'b010011000},{9'b011111001},{9'b000110000},{9'b001100000},{9'b111101100},{9'b010010110},{9'b100111110},{9'b110011111},{9'b000111011},{9'b011110111},{9'b001011001},{9'b110010101},{9'b101110100},{9'b101011110},{9'b000000101},{9'b111010111},{9'b010001000},{9'b100001110},{9'b110100111},{9'b010111010},{9'b011011101},{9'b101010100},{9'b000111001},{9'b011000110},{9'b101110011},{9'b001111010},{9'b101111110},{9'b110100101},{9'b110010101},{9'b000101000},{9'b011010111},{9'b101000100},{9'b100111101},{9'b010010011},{9'b001000011},{9'b101000110},{9'b111011101},{9'b110111101},{9'b001110011},{9'b110111100},{9'b001010111},{9'b101011011},{9'b111101001},{9'b011101011},{9'b111110111},{9'b000010001},{9'b111011010},{9'b000001110},{9'b110011001},{9'b001000110},{9'b101000101},{9'b110111010},{9'b000100101},{9'b011111111},{9'b010110011},{9'b010001111},{9'b100000101},{9'b111001101},{9'b111011110},{9'b011101010},{9'b010001001},{9'b010100111},{9'b101101010},{9'b011100110},{9'b000111000},{9'b101001001},{9'b000011100},{9'b011010100},{9'b011110010},{9'b110010111},{9'b000011100},{9'b101010101},{9'b010100100},{9'b000100000},{9'b011000010},{9'b011111011},{9'b111101000},{9'b001111010},{9'b100110010},{9'b101110101},{9'b111001110},{9'b001010010},{9'b011110100},{9'b010101101},{9'b000001011},{9'b001010010},{9'b001010011},{9'b011000010},{9'b111010001},{9'b001111011},{9'b101110110},{9'b110110001},{9'b111001001},{9'b110011011},{9'b111101010},{9'b110100111},{9'b101101010},{9'b110101001},{9'b111100011},{9'b110011100},{9'b001110011},{9'b100001101},{9'b001111001},{9'b010101000},{9'b011110010},{9'b010011110},{9'b010101000},{9'b000110101},{9'b111111011},{9'b110100000},{9'b111011101},{9'b001001010},{9'b111101101},{9'b011010111},{9'b011000110},{9'b010001000},{9'b011011100},{9'b111110001},{9'b111000110},{9'b010010000},{9'b010111010},{9'b001011110},{9'b011100011},{9'b110011101},{9'b001110100},{9'b100110110},{9'b111010100},{9'b010111000},{9'b011010001},{9'b110100110},{9'b111100011},{9'b001111111},{9'b110000101},{9'b111110011},{9'b010111100},{9'b001111100},{9'b111001001},{9'b001100111},{9'b000110101},{9'b111001000},{9'b000101011},{9'b000111110},{9'b011101100},{9'b100010011},{9'b011001010},{9'b100001110},{9'b001111110},{9'b111101110},{9'b011101111},{9'b001101010},{9'b111001111},{9'b111111100},{9'b011000111},{9'b001010011},{9'b111011101},{9'b011100011},{9'b100110000},{9'b111100111},{9'b001010110},{9'b011011010},{9'b111000000},{9'b111101110},{9'b100001101},{9'b101000100},{9'b101011101},{9'b111111100},{9'b010110111},{9'b110011100},{9'b101010110},{9'b110100010},{9'b111001011},{9'b011001010},{9'b010011110},{9'b101000001},{9'b111011101},{9'b001000010},{9'b110110100},{9'b110111011},{9'b011110010},{9'b111000101},{9'b111110011},{9'b111010001},{9'b100101001},{9'b000110100},{9'b111001101},{9'b000000110},{9'b010010000},{9'b000000101},{9'b100111000},{9'b111111010},{9'b101001101},{9'b000000000},{9'b101001111},{9'b001110000},{9'b111000110},{9'b010101011},{9'b000101011},{9'b011101111},{9'b011100011},{9'b011110000},{9'b011100111},{9'b100111010},{9'b100100000},{9'b101100001},{9'b101001010},{9'b010001000},{9'b010100100},{9'b011111010},{9'b101010000},{9'b111110110},{9'b011100101},{9'b011101011},{9'b000110011},{9'b001101111},{9'b010000010},{9'b010110101},{9'b000001111},{9'b010101111},{9'b010001100},{9'b111111110},{9'b011001011},{9'b000011101},{9'b010100111},{9'b100101101},{9'b010000101},{9'b011010000},{9'b011000100},{9'b111100011},{9'b000100010},{9'b101001111},{9'b011011001},{9'b110001001},{9'b010110000},{9'b010011111},{9'b101111010},{9'b101110100},{9'b000011001},{9'b000100101},{9'b010100001},{9'b110011001},{9'b000010011},{9'b001100001},{9'b101010111},{9'b111011111},{9'b110001001},{9'b110101111},{9'b000011111},{9'b101001100},{9'b101111011},{9'b111100101},{9'b100101110},{9'b110010100},{9'b011101101},{9'b111100100},{9'b000001111},{9'b001111000},{9'b111011110},{9'b001111100},{9'b111101111},{9'b110111100},{9'b000101011},{9'b001101101},{9'b011110000},{9'b000001010},{9'b100100100},{9'b110001001},{9'b001100110},{9'b001011100},{9'b111001100},{9'b001000111},{9'b010010111},{9'b011111111},{9'b011111000},{9'b001101111},{9'b101000010},{9'b110111010},{9'b010111111},{9'b001000011},{9'b111001111},{9'b001111001},{9'b000000111},{9'b110000101},{9'b011000001},{9'b111001001},{9'b100110111},{9'b100100100},{9'b100011110},{9'b101110111},{9'b111111010},{9'b101000110},{9'b100001010},{9'b000010100},{9'b010011111},{9'b110100000},{9'b100010110},{9'b001010010},{9'b101011001},{9'b000000101},{9'b011010111},{9'b110000000},{9'b101010111},{9'b110100110},{9'b111011010},{9'b011110011},{9'b010011011},{9'b110100111},{9'b001111100},{9'b011000011},{9'b110111111},{9'b111111010},{9'b010001001},{9'b100000001},{9'b101010101},{9'b101000100},{9'b011001001},{9'b110001011},{9'b101001001},{9'b011011111},{9'b010000110},{9'b110100101},{9'b110001111},{9'b111110011},{9'b000001111},{9'b010101101},{9'b001111011},{9'b100101100},{9'b010111110},{9'b001111010},{9'b001101000},{9'b100001100},{9'b000111110},{9'b001000100},{9'b100000111},{9'b111110111},{9'b001011010},{9'b001000001},{9'b111111011},{9'b001000100},{9'b111101100},{9'b100110010},{9'b011010111},{9'b001111010},{9'b111000000},{9'b000111100},{9'b111110110},{9'b000100101},{9'b010111001},{9'b001011011},{9'b100100001},{9'b011100011},{9'b000111100},{9'b111110111},{9'b111011010},{9'b011000100},{9'b000001111},{9'b110111001},{9'b001110011},{9'b100000100},{9'b010110001},{9'b111111011},{9'b110110011},{9'b101100111},{9'b011001100},{9'b111110110},{9'b100000111},{9'b101100100},{9'b110110110},{9'b100010011},{9'b111000011},{9'b011011110},{9'b110101010},{9'b001010101},{9'b000110000},{9'b111011011},{9'b001101000},{9'b111011011},{9'b111010111},{9'b101100101},{9'b110011000},{9'b001111011},{9'b110011010},{9'b110101111},{9'b111101010},{9'b100110001},{9'b100010101},{9'b010111000},{9'b100011001},{9'b011111110},{9'b101101001},{9'b000101100},{9'b111100001},{9'b001011000},{9'b011100110},{9'b100001000},{9'b100100010},{9'b000100010},{9'b110000000},{9'b110010001},{9'b011100001},{9'b111101000},{9'b100000101},{9'b110101001},{9'b010111100},{9'b111101000},{9'b000111101},{9'b010010100},{9'b010101011},{9'b100000110},{9'b100110000},{9'b100011111},{9'b111011101},{9'b101110010},{9'b000101000},{9'b000100110},{9'b000110110},{9'b011101110},{9'b101101000},{9'b010111010},{9'b010001111},{9'b010011101},{9'b011000011},{9'b100001100},{9'b001111101},{9'b111101001},{9'b111110111},{9'b010010101},{9'b111000001},{9'b111110110},{9'b110101111},{9'b101100100},{9'b110110110},{9'b001010011},{9'b011111011},{9'b011000111},{9'b000011100},{9'b111000111},{9'b010011101},{9'b011110110},{9'b111001111},{9'b110100001},{9'b110011110},{9'b111000101},{9'b110000010},{9'b010110001},{9'b010100010},{9'b110101111},{9'b100101100},{9'b110100101},{9'b010000001},{9'b011101001},{9'b000000011},{9'b011100110},{9'b001010111},{9'b110100110},{9'b000111011},{9'b110100101},{9'b010001010},{9'b010000101},{9'b101011111},{9'b001111001},{9'b110011011},{9'b110110110},{9'b001001110},{9'b100001001},{9'b001111011},{9'b101001110},{9'b111101110},{9'b100011011},{9'b010110111},{9'b100000111},{9'b011000000},{9'b001111101},{9'b110101110},{9'b110110000},{9'b010001001},{9'b011011010},{9'b000101100},{9'b101101110},{9'b101001110},{9'b011100010},{9'b111100111},{9'b100011010},{9'b000010010},{9'b101001110},{9'b100010100},{9'b111001100},{9'b100010011},{9'b010101110},{9'b011011000},{9'b011011111},{9'b011101101},{9'b011101111},{9'b010011010},{9'b001010101},{9'b111111110},{9'b111011001},{9'b110011001},{9'b111110000},{9'b001000101},{9'b011000111},{9'b100101010},{9'b111101011},{9'b000110001},{9'b101100011},{9'b101111101},{9'b001101010},{9'b101000101},{9'b110011001},{9'b101110001},{9'b100000100},{9'b111110010},{9'b110100010},{9'b010100000},{9'b111101110},{9'b000110101},{9'b010100101},{9'b010010101},{9'b110100101},{9'b000110001},{9'b101110100},{9'b011100110},{9'b100010010},{9'b001100110},{9'b001001010},{9'b111000001},{9'b000001010},{9'b000101000},{9'b110001010},{9'b010111001},{9'b101101101},{9'b100111101},{9'b100111000},{9'b001101101},{9'b011111100},{9'b010001110},{9'b101111000},{9'b110110001},{9'b100111101},{9'b100011111},{9'b001111010},{9'b010111000},{9'b001100111},{9'b001010001},{9'b111101011},{9'b111100111},{9'b100110010},{9'b010001110},{9'b111101011},{9'b011011000},{9'b111111101},{9'b010001000},{9'b110111101},{9'b010100110},{9'b100111010},{9'b111101100},{9'b110110000},{9'b110000111},{9'b001111101},{9'b110110000},{9'b000010011},{9'b001010011},{9'b111100011},{9'b101100010},{9'b101011011},{9'b110011110},{9'b011111010},{9'b011101101},{9'b101101111},{9'b101001011},{9'b100001011},{9'b111010101},{9'b001101110},{9'b101011011},{9'b011100011},{9'b101000000},{9'b111011101},{9'b000110011},{9'b000110001},{9'b111001110},{9'b101110111},{9'b010000100},{9'b011011010},{9'b001111100},{9'b000100110},{9'b100000000},{9'b111100001},{9'b000101101},{9'b011100100},{9'b100111100},{9'b111111111},{9'b101111111},{9'b001000101},{9'b011000011},{9'b101010011},{9'b011111110},{9'b010011111},{9'b110011111},{9'b010101101},{9'b010001010},{9'b100110001},{9'b110110111},{9'b101110111},{9'b010001111},{9'b111011011},{9'b100100011},{9'b101100101},{9'b000011100},{9'b111110111},{9'b010101001},{9'b110100110},{9'b101001111},{9'b111011001},{9'b101100001},{9'b100001110},{9'b001101101},{9'b111010100},{9'b000100011},{9'b010000110},{9'b111101101},{9'b111111100},{9'b010111111},{9'b101110101},{9'b110011110},{9'b011111011},{9'b010001101},{9'b111000110},{9'b101111111},{9'b011001111},{9'b000110010},{9'b011111011},{9'b110101000},{9'b111101001},{9'b111011101},{9'b101100001},{9'b110010010},{9'b110111001},{9'b110001010},{9'b110101100},{9'b100101100},{9'b000101011},{9'b011110000},{9'b001100000},{9'b011000110},{9'b101010100},{9'b110000100},{9'b011011000},{9'b111010101},{9'b011010101},{9'b000011010},{9'b011110111},{9'b011111010},{9'b101010101},{9'b000101100},{9'b001101000},{9'b111111100},{9'b000111111},{9'b100011001},{9'b110110101},{9'b010010101},{9'b101100100},{9'b100001100},{9'b011110000},{9'b101011110},{9'b001101100},{9'b111010111},{9'b111010010},{9'b101110001},{9'b000111111},{9'b111010011},{9'b101011010},{9'b001011110},{9'b110011010},{9'b111010111},{9'b101001111},{9'b111001101},{9'b001110101},{9'b001011110},{9'b011110001},{9'b110110111},{9'b001010010},{9'b101111101},{9'b000110001},{9'b111100100},{9'b101010000},{9'b000010111},{9'b101100111},{9'b010010110},{9'b111010001},{9'b101001110},{9'b110101101},{9'b010000100},{9'b110111000},{9'b010010101},{9'b101000001},{9'b001010111},{9'b001001000},{9'b000110000},{9'b010101110},{9'b110111001},{9'b111010001},{9'b010110111},{9'b100011000},{9'b110110111},{9'b110111101},{9'b110011111},{9'b010010011},{9'b000001001},{9'b001011110},{9'b011010011},{9'b000100110},{9'b110101101},{9'b010110001},{9'b001000010},{9'b111101111},{9'b010000010},{9'b101011111},{9'b001111100},{9'b001101110},{9'b111111010},{9'b100011001},{9'b010110001},{9'b101101001},{9'b001110111},{9'b111010011},{9'b110110111},{9'b100101010},{9'b010110010},{9'b011111101},{9'b000100010},{9'b110010001},{9'b110011011},{9'b011101010},{9'b100101010},{9'b100000000},{9'b100001100},{9'b011010101},{9'b110011011},{9'b011110101},{9'b100101101}};
assign weight_o_4 = {{576'b000100110110111011110100011100100100101101011000101001000110001110110011001011001111011101110010100111110101101010100110011000101001001100101100100011010100001011001111000111001000011101000001010010011101011110111000010101000000010010001101001111001010100101010110111111110111011110010010110110001101011101110111011011001011010000101001111111011110101011001011010001100101011101100100101000011101101101100000001001101000111110111111001101111111000010010111001011111010110101111010100011111100111100000100011001111011001101101111101101111000011010011101010111001001011011000010},{576'b010001101000000001010111100110111101100011111001110100000111111010001001001111001011011101011001010001101011110100001100111100101111001100001100111010000110011000001110100001100000110010010001011101111011111110111100010111101010101110101111100111011011000100110101100111110010011000100110110110100100000001100110111000010011001001010111101000111001111011010100111101010111001011001110010001011110101001111100101011110100100011010011011001111111110110101010010101101100010011110011110010000110100100000000000001110000011100111001011001101000101011001111011110110110010001000010},{576'b011011101100110111111100011000000000100010000010100110111011010100111101101110100111011000000110110100110111001011100110001000110111000111010111111101110001010011010100010101100110011110001010110000101000000001010101110000010110000001100100100110110011010000000000110000010111001010111101000110001100011011111111001111001011011100100100101011000101001010111011010011001000100111001011000101011011101001100100111100101000101100101010100010001100010110000011111011010011100110001110000101111011110101001100001110100011011101111111011011111000101011011010010101101011011001000101},{576'b001010111100011111010001001000101100000100001010100101100110000100011011011011101001011111101010110111110110010101100000010001101010101000111111111011111000011011001100010111001001011001000010110111001010010110001000010101000010010010001010100010011011110100010011101110100010011001110000110001111011101000100000111101010111001111111110001001010111101111001011010010010110001101001110100010111101111101011100011001100001010011101101011111101011111011100001110101110011000110001010100111011100110010111111101010100100100111010111001000000000110000000101101010000111111010110010},{576'b110010000101011010101011000100011011010010011100100110101001000100000011111110100010010101101000110111111010000001100010000010000110110011001001111110001010100100000101100001101001111011110101000000111111001100110011101010101101110111001110101111111110011011011000000101101000101100001011001101001111010011010011101110001010011000010001101100111001101000111001111101101101110110110010110010001101010110111000010101000010110100001101101111101111010010000011001110000100011111011010110010111111101101111100010100101101001011010110100010101101101010011101010111001010011000001110},{576'b100000101101110110010011110011000000011010101001010111001100001010111100001011011010010101101010101010110001110100110100010000110000010001001001111110010010011010011001000000101111011111100100000010011101101010100000001001000000010010101000011110101010100001000101110011011101000010010000110101001000011000001111101000001110110100011101101110000000111111001010111111110111110010111010000000001100011101010011011011110101110010110001011101101010111001001010010100101011011000001001110101010111000101110010010010100000000110111100011000010010011000001111101010110010110001001010},{576'b110101101000001001010011110111111111100011111011011110110110000010111100001011001111110101110101001010101111111110001000011110100010001101011011011101111000111010011000110110100111011100101110111010000101001001011000111001010010100010001111011111111011110010010010011100001010010111101010000010110000100010101111011000101111111100101100111001010111101010001011010111110000010101000010101010110111110110110100011110011000101100101001000011000100001100010111101111010011111100111110010111110100000111100100010011111100101101110111001100010010110000000111111010010110111010001011},{576'b110101001100011010011000011100111000010111001101101110001011110011111111111011110101110011110110011101110111110110000000010011110001001001110111111011111101101110010011010111101010001101001111100110000111001010101111110100001111011101011100101110111101001100111001110011011011000000001100010001001000100000101100100100000111111001011011011111100011111111001000101101101011010000111011110000111110101001101100111010101100111010011000001111111010110110100101111011011111111101100100010010001011011001110100001101011001010101111001101011011111111000110110100111101010110001011111},{576'b111110100100011100001111000110101111111000111100101100101100101101100010000100100100011111011011111100000111001101011011001110111111100001001000010000110001000000100101001111101010110001100001101110010000111110101100011010001010100010001100101111001001010100101001111011010010000101100000010010101000010010101111101010010101000111011111001011100010111101000111011100010010011001001011110010000101101011001011100101111101010001110101110100101111101111110110111110110111110001101101110110001011001111010011001110011000100110110110101001010100111000001010000111001001011001000111},{576'b100101101011000100011110101111110111101111110011101011100101101100110001110011011111000101101000010010000000101001001011100000010011001110010110001011111001101001110010010000010010011101001111011110101100111011101011101001111101100001110110001100100100101000111011000000000000110111110011011010100100110010100011001001101000001001011000011101111110111111101001101101100111001100111000110001000010111010011101110100011011011100001100101110101110010110010101101111100100111010010010001101110101011100101000010001011111011101111101010010100010110000101011101000110110110010111010},{576'b000111000001111101101110101111111111011001110101101101000100101100110001100101100110111000000010010000110100001101100011010101111001110110111110110010101101011011011100011110011010001001001110011110000101111100001111001111101111011000110001101101111101101111001101001011111011100101010000100010010100110010111100111001110010010111110110111001001101001010000001010010110111001001100111011100101101111001101111110110111111000001011001001100110010111110000110010111100101100111001101011101011011000101111000011110111011100101001111111110010110100010001000100011100001111111111011},{576'b001010001000001000000011001001000001011110101001010011000111100100101000110000101001000111000010100001000000010010011010111000000011011111111011001011110010101110010011100100011110001101111111011100001110000111110000001001100100100000000110111011111010010010110101010011110111111000001001100110001000011000110111101111010100111000001010110000001001000110010100001000001101100110011001100010110001000010000011000011011100100110101110011111111011100110100101011011011010000101001000000010000100111010011100111001001011001101110001011101100011111110111001100100111110111101101011},{576'b111100100101101011111111110011111101010000110110101100111110101110100110001010010101001000100100011011011010011100111100110110101000010100111101101011111011011010110111110011011010011001011111001101001111111111111101001000110100100001010011011001110110010011101001110101100011000101101100010000001010101011111001101111010011000011101111101100000010000001001000000010101001101010100100111011110011111000001100011101100110011000110100001010001101000101110010110101000001010000100011010101001011100111011000000100100000001010010000010000111011101101111011101100110010001001001110},{576'b111001010111110101110110111111011001111110011011011001010101111101110011000100000000011111011101111110001111011000011011000110111111110100101110101001010111001101100010000011001010110111010011011100101101001101101111000111111101100011010000001001110001101110100101010010101011000101001000000001001000100000011101101110001010100111101011111000111010110001100101000001111110010101100101100111000001101010101111111100111111011000011100101111001101000110001101011101111010110101101000100000110001110110001100010011110111011110110000001011100011111101110110101100111100010001001111},{576'b101001110101010000001001011011000010001110101011011011000101101111111101101010101011110001001000100000001100100010111000101001010111100101100010000011001111111100110110011100010010101110001101010110000101001011001101111100011111011010010001101001111101111111101000011000101000110001110000101000110010100000100011110111011010100100101000001100010010101010001100101011010001111011000000010010001100000100101001001011110110000100110010001100010000100111101001000010100010110001101101110000101001001011000011100111000111001101011001001101000110111001000110100010001011011110010000},{576'b111010010110100010101100011110010110011110000100101011001101111111101010110000100000101110010001110100100111000010100001110110111101101010000000011000010001111111111000101100010110001100101011101010000001010110001111010111000010100110001100001011000111101100101001000011100010000101000000000000001000100000111110111110010010100110000111101000010001100011000011100010000001111010111001010110011101111100101010001111010101000000110000001000100001110101111011110010100000100111010101010101010010000010110001110110010111101110010011000010000111010111001001101100100100000110111000},{576'b100001000011101100101111110011100001011111111101101101101101011010010110000100010100111010111111011000111011001100100011001111110010000110011111001110010000101010001000100010000001110010110001010111101101001110101110010111111111000011110001100100010011111101110010110111100110101000010011110101000111000000010001100010110010101011010110001010010110101110001001100010000101111000101111111111100110000111110101001110101000100000000010010001010010000010101000011001001001011101010000110001110111111010110000110000001101010011111111110011101111111101110110011101111010001011010100},{576'b001011001111100101001010001111000010001110110011000011010000101001011000110001001010111000110001010001000011000000000000100000010001010010010110000010101000110110010110110000011110001001111101110111000111111011001111110101010111011001110111101000100101111101111010010010101000011000010101111101101011000000100001100110011010000100101010001101011101100010011001110011101001110011001110101101011111101011110111110011101001000011111101111101110111101111111010010100100000001001011001110100011110100000100011100110101010110101111010001000111111111100110001111001111000111101101010},{576'b011010011100101110101001001000101100100010001000000011111011000101001101101110000111100100100110000011111110010101001111011110100010101110001110001000100000001011000100000011001011001111000100010101001011100111111110001011110111101011110011011001010111111001110001100011010011100100101010100010000000011001011101001000000010100111001011001010010110101010001000100100000101011110000001010010110000100010000001010100010100011100100000010110111000100000101010100001110010001000101000001010001000000000011111001010011011001101101101001101011000001000001010010011001111110011001010},{576'b000001001111010111000111001110010110100110010111001001110011111111101011010010101000000001111001111000100000000010001001100100010010000011100101001010000110111010101001101000010010111010011100100011000111110100001110101101010011011011110111101011000101111101010100111111110111110000011111110111101001000001110011011011011110111100001010010101111110011010011100111010111010011111011000000101011000011100111001000010101000110010001000011111001110000110111011000011000000100000110100111001111010000100101000100100110011011110100100011110000000011110001001011110110101111100101010},{576'b010100001111000101001011101111111111101001110111101100110111111111111101011100111010111100111101101000111001101110100101000011110010101010000000100000010111100111111001100000000001001100100011100010010000010010001101011110010010011110001000000011001000101101011000110111110110101000100101110100000101000001010000011110111010110100101110101100010100000010001000100010101101111110100000001100011110000110100101001011000000101010010100101001011011110110001000000000101000010101110000011001110000110010101110110101111101010100111101100111101010111000010110111111111010010001011101},{576'b000111101011000101001110011111110111001011110001001001000001101110101101001100001000110001111100001100111111110110100101000110110010101100000110001001010100101010001101000010001001111010000100010101011110110101101100011100110101111001010001111000001100100101010111100111110010010110000110110011100111000001100110011001000011010110011111101010000000001001010110011011001111010011001101010011000101010001011100010110010110000011111100001110111010100110000011100110001101011111001001110110110110011001110001011000100011010010101110111010111100011111001011011001000111101101100010},{576'b001101010101110110001001011011000100111010101100001011001001100001010111001111111100011001000110110110000100000110100101110100000011110111001111110000010100001101011110011001001111000011000100111101001010101001010111100101111110011100011110010000010111000001010001101111000100111011000010010101001111001010100011111011000000101010110010111010111011011001010110010101101000010011000010100100011110101011101101010000011111001100010110100001011111001101010101111011010100110000110001010111100111010101101001000000011010000100011010110000110101100100000000110011010101010000101010},{576'b111110110111011100001111010110111111100011001010011111110101101100000111111001011011110011100111010111100000001101101110100011000001000110101101000001100110100001000111011110011110001101001101111000000010101011001011100110101101000000000110000001001100010000110101111011011010111000100010010101110011000111110000010000011100110101011100011101100101000001010101011111110101010000011010000001011011101101010111011011011101001001100101110101000111110110000001000110100110011111010100000000011110111001111001001110110011000110011111101010100001011011011100011101100011010011010001},{576'b011101011110110110111100101100111101111001100010111011011100110111000110001100000001110011011100000110101001101111101111101111101011110111101111010001100001101001110110011101001111001001000100011101011100110000101100001101101101111000010001011001001100011101110111101010000100100001100101110111100100001001101111110010010011010111001110110001100101001001010100011111000111000001000101001010011101011100101010000101101111100110001110000011111101101101010110111001111111100010110111110111100000000101100110000011010011011110111110001011010111011111011110100000100110011101101100},{576'b110100000001110100111100011111010100011010111001100011111011100000010011111000010111010111111001110111101101110001110110111000000100100011011000000110000110110100010100101110010110101110111100101010011101011011000111000110001000000110011100000101001111011001010101101011000000100001110001010111110111000101101011011011100010100000101110000000101110011101110001110001010001001000001110000101111101111101100100110110101100110011000101001111101110101010101010000101101110011111010111101000111010110000010100011100101000100100011010010101111000011010000011101011000011010001111010},{576'b010010001100110110101000001101001100110010000110000011001110010011010100101110100001001111000100100010111100111111010111111111101111000111011111101000111001001101011110111011000001010011001010110110011011101110111000111011000001010111100011010010111011110000010111000111100000101001100110010110100101000011100011111001111010101110111100010101100100000001101010011100110101100100110011010010010101000110111000001001010011011010001000101111111000100110101110001001101111111111100010110100110100111001010100110001101101101100000010110000100101000110110111011111001011100110010000},{576'b110000000101000001010111111111000001100010011111010000010010111001000011111110000011010100100101010101100011000111111010001010000100001110111000001110000110000100011010111000100110111100101101100011010000100001010111100011011010101110001100101011100111100000010111101111111101001110000110100101110110111011010011011100100111011111111001011101000111011101110111001100010100011010100110110010000001001010110111100111011010011110001110010011111111000000010001110111100010110001000000000111111110100011111111110111000111011110011110111001101000001111011100010001101111010111000010},{576'b000101111110010111011100111001110101110001111011111010111000110101110101111011010101101010110110010111100111111111101011010010010100000100110000000111000110110101001110110110001010101110101000000000110110011000101000100100111011111101001100001011101100011101111011111001010000110001011111011110000111001010100000100010010011010110011110001011100101111101110000111100010110001100001111011110011100010110111111010010110011010001010001001100001000110110011101011011010101010011101000010111101011101100000110001001000011110011000010110011101001100100110000011001100111100100101111},{576'b110100110111010100101110100111111110101100111010001000110101100101011110011111101100101001011001100001011111101001100001110001011101111000100010111101110101001110110001011100011111010101001111011111111100110011011100000110110111010001110001111000001100010000011000011000000101110110011110001000001101010010011011110000110111011000001110101110001100101000111000110100110111101011111100100000011101011110110100100000001111011010000100000111101111011110110010111101101110010111100010000000111100100010110110011001100111101111000101000011000111100100111100011110110110011100000101},{576'b010010000100001011000011100011110001101101101101110100001110111100010010011000000111110101001111100001001011001010111111100100110111110111111110101111000010010001011110001100111110110011110001011110111010001011001100011010010011000101100010111000111000110111100011110100111011100010000100100011011000100011111111111001000011100011000011000000000001111000110111001001000011101111000011011101111110001001001100100010110111101011111001011010101100110111110000101011101000110010110011010110000110010101101001010011101001011100001011011101111101110110011001101011100101001100101110},{576'b111110011101110101101110000011100101000001100100001100101100010101111111110111010000110001011001011111000111001101101010110000011000101000101010100110001111010100101001100010110000101100101011011111001100010011000100100110110011110101110101111100001100110101111101111101010000010000111110011101101110000111101100000011110111101110010101000011000101100101100100000100110010101110011001010110101100100001000100000111110011010001110000001000001100111111111101110111111011111110000110110111100100110000001100111101000111011110111111011011000011110101011100011100110001001011010000},{576'b011000110101001000110100111011011101000011010001000000110110001111001100001110101011110111011100100000111001100000111011001110111111110101111111111111100101110000000010011110110000000001110010100000000000100000011000011011000011001111110001110010101011110110000010011010111111011110100110000001111110110011110010110001100111011111101010001011100110000110111011100100110110101100101011111100100110101101110001100001101101100110001000011111110110101011111111110011100110111001001111110110001101001100110001110001011000000001100000101100111010001010001111110011100001010100101000},{576'b100100100101001011110011010010010000000111101111010000110011011011110101100011111111100110100110110101101011110011111110111001001011011000011000100110101101001110011001110101111111011101101110000011001000100010011011000001011001010000110001001100000100001101001100000010101110100101111000111110001000111110111001101010100101100111011111010010100101100101010000011100011100000010001011001111111111100001011111001101110110111111110011011000110100001101110111101011010001110001101001100111101000100101101111101111010011010111111111101111001000011011001111100011000010111011100010},{576'b110010000010000011101001100100110011011100001000100010111100110110000010001011110101011111110101110000011011110101101011001010110111111010100000001001000010001101100111001100110100101100101010010101100000110000111010110001011001100110100011111010110011111000101010111000110111011111101111001000000101110000011100000001110001000011010011111000111000111101011001010011011011001001101111111110000111001000001100000111110011101111110101110111011000000110000010010010001001011111101100100011011100110000111110001101101001110010111110001111100001011110110001100110111111001101011001},{576'b100110011100111010100111000110010001000101000100101100000100111101011111101101010000110001111100011110100101001110100100100011010111101011100101010011000001111100110010001101011110111100001011100000100100110110110001111001000010100000011001111010101010101011111000110011010111110000101100110011101001110000111100111100101010101010000000100000000111100100110000010100011000010110000011011010100001000000000010011111010101000001010001100100110000011111101010110000101000000100100001000000000100000010010000100011001011010101111101001110011110011000001110011111101110110011110100},{576'b000001001100000011100001111000110001100100001001000111000110111011101011001100101110001111111001100000111000101010000101101001100010000001010010111000011110001100100011100010100010001111101110111010100100001010000101110110010011000101001000100100111000111101101010110001001000101011001001000101000111000110011000110011000000000101000100001101010110100110001000100010110001100000100110101110110000101010111001110100101011111011101100110011001111100111101100011001011011100110001100111111000110111000101110001010011010010001110111001111011010101110001000010011010111010001101110},{576'b001011001100011010101000011110011011100000110001010000010000011100001010110000001010100101100001000000010000100000010001101011111010101000000000101000010111100110101001100010100001111000100110110111111111100101000110100101100011011100110010111000010101100110101010000100101100110101111001101100010100100010000011100011111000010101110101011110010010111010001111100010100111111000110101100010001100000011110000111010010011110101100001010100110000001101111000111001000011100001111011000010001101100100101101001011111010010001111111111110010100101111101010100010010110111001101011},{576'b011101111100111011111001111000111000100110101100001110000010001001010110011000010011111010000110110001000111010010110000110011001111111000001001000011100101110101110100010100101001000010010001111010010000111010000101011110000010001001001100100110010001001000111000110001011000100011101001011110010100010110010000110011110100100011010101100010000111110100110000011110010000010100011011111010111001100110000100011111010111010000010010100001011001100101101010110001011010000000100001000100010101100000011110100011111101011100101111011110101010011001011100011001001111011011001000},{576'b010111111001111101011100011111110011010000110011111111101001000101101011000000101010001101101001101000011000100000010001001111111110101101001010001001101111000011100011000011111010011101010110101100110111000110110101011011100100111100011000001011111010100011110011011010101011100001110100100101110000101111001111000110100011001111110111111110011010011010011001011110010011111110101110111001111011001011000100011110111010000110010010100000110011011100010111111111010111110011101111100011111010011101101110011100001011000111100101101011010110101000001010000110000000111110100100},{576'b000000101100011111110001001010001000100001001101011111110010110011100110011100101111001110000010100010100111110001000111011011110001011110111101011110111100011000011111111011001111111011001000111111100111100001011101110110101111101110011110100001111010001011101000000001001000000101101001001000000000010010010000100001001010111000101010100001001111000011100010101111101010001110000010101010111101101100000100110110010011000100010011100000011000100100011111100101010100111000111111011010111011101100100011001010110111011100101000000111001100011010011110011010111110110100011011},{576'b000101011110110101111100000011100100111010101111011011101111000100101001011001100010000101101001101000000100000000010000101001110000100000011010111011001010000010010110101010111001110011000010100111101111100011010010001111110111000111110011110001110010001011101011000100001010110011001001100010010101101010001110000100111110011101000110011101001110101110001000110011010001011001101110111010000000011010100001100010010010100001000100000110111010010101001000111110011011100001111111001010110111010100000100001000111001011101011101011110111110011010001111100011000111111010101100},{576'b101010101111000111010101000010100100001110011010111001110011101010101000010000101010001110001001110100100000110010010000100011101111111111011011010011101101010101110110011100101000001110011001001010001101001010000000011110011111000001011001100000000000001110101011010011101000011101011000001001110010110110000001100100100011001100100111001111011110111011001110011011001011111011010000011100101110010101001100001011000110111001110010001011100100000101110111101011110100110011101100010011100111000111101011000011010111111111101101000011001111011001111110011101111011111000000101},{576'b110011011001010111001001010110111011100010101101010011111010111001111111110111010111110000101110111111100111111110111110010100000011000111001101010010110010000001101110011001010100010001001011101100110111000101001110001011000010101001111110101101110000001101110111111011010011110000101100010001100101001010010110100001010111100111001101010001000110010001101110011111011100100000000001110001111111001110110001101011011001111100010010100001101111111001110111101010010011110011111011010101100101001110101111110111010001100011101100100000000010000101011110011000010000000011000111},{576'b011111111100111100001110011010011101110001110001111001000000011111111011011101010100010111101110101010101011101010001100001000011111110001101101110010000010010110111101010011000101010001010110111111011110100101110001110110101100000001000111001001110011000010010100111001010100100000110111111011100100010100101000011000010111011110111101011111001000111000001110110110101010111011011101010100101010011110101011101001110111111101110101100000000000111011111011010101110100010110101110100001101001100010000110000001111101110111110101110000110111110010010111101110001010111010111100},{576'b011000101010001111110110100101011001011100000011111100111101111010101000001110101011101101010101001110111000110101111110011111100111111111001101000011001011001001111000010100111111000000011111011110101110010101101110101111101110111101010111001011110100100101000011001100100111010011011001100101001001101010101111101110000111010111101101010011000010101001101110010111101111111001000101101101101110001001000101100010001010001111001110000000011010000101110010011001010100101010111110111010111011111000001110000010010111010111101101010011001010010001101100010101111011100001000011},{576'b000011101101111011001000111100110110110001100101011100001110001101110010111001001110100100111011111010110000111000100100001000110111010011101001110010011011110101101110000001010010010101011000000000110101001101111110110111011010000110011010101001111011110001010001010110010000110101101000010111000111111000110110011111111100100000110010010100010000110010100001101011100000111110111000000011111111111001011100111011000001010001111101110101100001011000100011011101010110101111011001110000111110101000100111000011010100100011011110100111000001111101010110001101010100001101011100},{576'b000101010110100101011100011111010110110101111101011111110111111110001111000110000111011101001000100000111100111010010100001101100010011100011010001101111111000010011111111101111111000101111110100011001101010011000111001101000101111100110001010000001010011001110111111110010011110011011101110101111011001010101111011110000111010111101111010101000110010001001100011010010100000111000001011101110010100000111100010111011101011100010010101000111111100001110001100011010100110000100110011111000101011111100010010010010011011100111011010100111100101000000001101010101011001100111101},{576'b110010110111001011000011111111001010001111101100000011111010001101010110111011011000100010110011011111110011110010100001010011100101000110010010101000000000110101010100010000111100000000000101110000010011001000011011110010011001100110100100100011101011100010000011011100110001010011101100101000101001101010101111001101010111001100110001011111001111111010010110010100101010111101011101000000000011001011010111100100011001001111000010111001010011111001110011101110110111111010100010010101101101000011000001100111010011110101110001011001011110100010101011111110101110111100111100},{576'b000010000001101010110011000011011001000110010001010101111011111001110111111111010111111011111101110111100001001011101111110111010011011111001111000011000010000101001100011001010111000001000101010000001110010100001000001101110110100101010110000111100100100101110011011101010111110111001110101000101001101010001111001101011100101100100011010100001100110011000110100010101010111110111001000110011110110011001010001001100110110001110001010000001101010111111010011001010000110010111000000001100101101000001111000000010111001101101111000111001111110000101000010110110100001100001101},{576'b011101111110010101111100110001100010010001111010100101110000010100000010101100001000100100101100010101110010010101101010110010101111111101001101000111101010111110111110101111110110111000011100001110100100110001010111000111100010100111111011011001110001000111000011000100010001111011101011000110111101100110001110000110110111011111101101011011001100011101011100010110110110011010010100110110101110110101001100001001100010111001111101001110001000011111010000101110001011010110001010010101111011010101111001100011001111111100101100001011001101110011110100100110101000111110010101},{576'b001101011111110100001100001011010110011000110000011000001100101101110111111111110110111011001011011111100111000111100010110011101011101100110011011011011110001010001010110111101001110010100111001101100101110110001100100000000010110001101101001111000100001110000000000111100101101110101100010000010110110000000101001011110000000011100101100000000011100100001101001100001101111010000001111110110000000100111011110111111000110011011010100011111001010000110100011011011100100100101111111011111010010000101011011010110011011101110101010011011010001001000110110111000011110110110101},{576'b000110101111100001001011101101101010011100111101011000001001110101110001111011111010101011010011111101000100000011101011111010001111110100011111010101100101111111011001011110011111001000101010011111111110110101101100110101101101010000011011101111101001010110110011010001010100101101111001001000001001101000010110001100011010001100010010111101111100000010000000100011101000011110110100111111110110010100011100000000100010110001111110101111101000010010110010001000110100010111111010001010100100110000010011100000110001101100100101000010101111110100100000110110101001111000110001},{576'b011110110110010100011100100011110011111001011101110111000101010100111101111011010100111000011111111101110011100111100010111000111000100100100101010010001111100000100010000110100000010111000011000000110000000100101110101011000010001010111010011101110001101110000011001100101111011111011101100100011100101011010111001111000111111111111101110111100001111110010100111101111011000001110011100000000010001010011111110100011100011100000111110010010100101111010111011110000011100010000010001101100011101111101010100011111111011111110111011111011110111110001000001110110000111110010011},{576'b001001000000101011011011001110111110010100100001001000110110100001110110011110010101111000011100111101101011001111101111100100111000011111011001001101001100001000001101111010111101000100100110011101111001100000111100010101111111001110110010110011110011111000000000111111001100001000101001010001110011000111101010110010110111011101110011010111100101111010100001100110101010011100110001110111011100110010100100011011100111100001100101010010000000111111111011001000100111001011011000110000011000001010001111101101000111111111100101001111000100111000001000010110100001111110000001},{576'b101100100000001001010111111100000010000011011010100100010011011100000000011100011110001110101110000000110110110011011101110100101011100001101100110000110010001101100101001100000011100101001001110100101000111001000000100010100101010101010011100000001100111110001000100000101101001101011000110101110000000110100011111010101100001100101010010100011110100000001011111110101010111100111000011101110010001101101010110011011000100100001010110011010001110110010111001110100111111111011011110110101111000001110011111111100111111110001111011011011100101001110100010110111100011010011101},{576'b100100100001001101110001101010001000101111001110010001010011010100000100000110101111010011100101100101110110000101100011101111100111001111101110001111000101110100000100101100110010011100110101011101111101111101101100010001110111110001111011110100001000010100101001011001010000101001011001000010000001110000010110010100011001101100100110010001011100101010001011110011100000111110100101100010010000101010110001111001000000100101001111000011011011010000110000111111111100011000100011011101110010000100100000111000111000101100010010000111111110000000101000100011011001110010010111},{576'b110011110001111001110100111010000000100100001111000001010011011110011111011101110111100111000010100010111000111000001110101101101010010001001110101100010110000001111111011101000010100011001010101100110001111001111101111010101110100010001110000111101011100110100011000100000111001111101011100010001110101110010100001001101110101000000010100110011101101001100000100100111001111000011001111111110001111100000111111010111110000001001100100100001001010010001110010101011011100110010111001011000101111101001100100101110011010100001010010101101001000011111101100001101111101011101000},{576'b111110110011001100100111110111000100011000001110100001011001010000111101111011010111010000010101011001100011101101100010000000001011011001101100111111001101111011111110001111111110101001110000100010110001010110110011011010000000101010101100100111101000001110001110011101011011100011000110001111100101111111011100000011001010010100110011111101111110100011001001010011001001101011111110010010001100100000000001001000010000010101110001001100001000000111111011000001110010111111101011110010001000110010011111101101100000110111111100011111100001110111100110011010100110000001100000},{576'b100011010001101000110100101010100000111011101001000110101111101100010010110101100111110010011011100001110101101100001110110110010111110111001111011011100111010101010100001010000010001101100000111101000110101001111110100101110101010100111110001100110110101001010011111100010110011111011110110101110101111010000111101101000000101000110011000001111110100100000000110101001001010000000101101010110001111010100111110000001000000001001100100101011111011010011111000001000001110111001010101010101010111001001100101000101010100100001110100010010111100000101000100011010001110110000011},{576'b110010110001000010010111111010000000101111001110100101000011010111001110010001001011110011101110101010100000110100011110100001110101011011101101110000010001011001110111001100100110001011001100101010010000110100001001111110000010100001111101110100010000000100101001010111101111010111101000110011111000101100001101001101101010001100011010100101111111000011000001100011001011000100110110111000100010001011110101111010100101001110011010001011101011111011100011000110101001000111110000111010111000100110111000011010100101011111100101001010110001011011111111100100100110111000101001},{576'b101011010000011100100111011000011000101100001100100100000001011000111101010110100101011000010001111000000111100010110000011000001010001111101010001111010111101000100011100011101000111000110101101101110110110011111100111001101101111110111111011011100111111011010111111100000111111111111111110101111001001011101110001110010111000111100110110000100001010001110101111100000010000011101001100000110011001000100111111110001100000010001110100101111011010110000100111011011111000111101110010111110100110100001101110011101011000100111010001001111100000111000000010011001001011110110110},{576'b101010100001001010010011110100101000100011001110100101011001010110101011000010100000110001111001110000001100100000010101001101111000000000000001101110111011010000101111000011010010101001001011001010011100110001101100001111010110010001111010001000000100000011101100000011010110100001001010111111000000110101011010111000000010100100001110000000100010000101001100101000010010100101101011101000010001101001011110011100001101000111001100000010010110001100111101000111110010011011111000010000000101111010000101100101011011110101111111011110100101001011110100100010111010101011110000},{576'b101111110101111100011010110101101110111000001110111011111001000010101101000110101111000011111000101001001110110100011000101000000101010101101000111110111011011001011111111000110110110011101010001111011011101001110111011000010100001101000000101001011001011011011111111101010010000011000110110111000101111001011110110011000100101000000001000001010110110110010100001110001001000000000001101010010001111000010111111010001000100010001100100110001001011110100001000111101011001111100000000010010000110110110001111101100110010011001101110000000001010101110111001100000110001111001001}};
assign weight_o_5 = {{64'b1101110010010001010011010101001110100010110010011001111000111101},{64'b0011001111000100101000110111111000010110101001110000011010011010},{64'b1011000101111011010100101001010001100011000111000010110110100011},{64'b0000011111110110001110110111111000100101101001101001100110111001},{64'b0010101100100100011010001101000011110011000110101100111000101100},{64'b0101001111011000111000100011110011000110010100000111101000011001},{64'b0010110011001111001101100101000011101111000101101001101001001011},{64'b0011001000100010010001010110001111001011010100100101100011110111},{64'b0001011100101001110001100111001111010101101101000110010001100000},{64'b1011010100111101100101010100001001101010010101101110100001101101}};

// assign threshold
assign threshold_o_0 = {4'd4, 4'd2, 4'd1, 4'd3, 4'd0, 4'd3, 4'd0, 4'd2, 4'd0, 4'd1, 4'd3, 4'd2, 4'd1, 4'd0, 4'd3, 4'd1, 4'd2, 4'd0, 4'd2, 4'd3, 4'd4, 4'd3, 4'd3, 4'd1, 4'd2, 4'd1, 4'd2, 4'd2, 4'd2, 4'd3, 4'd3, 4'd1};
assign threshold_o_1 = {9'd369, 9'd386, 9'd189, 9'd236, 9'd230, 9'd276, 9'd742, 9'd219, 9'd570, 9'd404, 9'd236, 9'd279, 9'd140, 9'd937, 9'd147, 9'd68, 9'd281, 9'd390, 9'd301, 9'd651, 9'd158, 9'd250, 9'd423, 9'd139, 9'd163, 9'd191, 9'd86, 9'd59, 9'd98, 9'd37, 9'd35, 9'd248, 9'd425, 9'd420, 9'd403, 9'd199, 9'd503, 9'd248, 9'd31, 9'd273, 9'd89, 9'd399, 9'd79, 9'd220, 9'd241, 9'd163, 9'd271, 9'd465, 9'd390, 9'd138, 9'd106, 9'd129, 9'd412, 9'd242, 9'd583, 9'd283, 9'd120, 9'd213, 9'd465, 9'd348, 9'd291, 9'd99, 9'd256, 9'd202};
assign threshold_o_2 = {10'd300, 10'd676, 10'd508, 10'd227, 10'd207, 10'd206, 10'd499, 10'd80, 10'd605, 10'd450, 10'd988, 10'd70, 10'd641, 10'd375, 10'd1248, 10'd221, 10'd235, 10'd261, 10'd659, 10'd469, 10'd706, 10'd581, 10'd42, 10'd146, 10'd101, 10'd699, 10'd402, 10'd324, 10'd115, 10'd103, 10'd151, 10'd129, 10'd1058, 10'd286, 10'd829, 10'd103, 10'd1107, 10'd220, 10'd46, 10'd60, 10'd481, 10'd543, 10'd435, 10'd193, 10'd498, 10'd218, 10'd329, 10'd85, 10'd544, 10'd194, 10'd109, 10'd761, 10'd385, 10'd290, 10'd317, 10'd1792, 10'd299, 10'd591, 10'd202, 10'd125, 10'd463, 10'd168, 10'd278, 10'd236};
assign threshold_o_4 = {11'd1029, 11'd191, 11'd677, 11'd471, 11'd2234, 11'd124, 11'd746, 11'd53, 11'd840, 11'd8, 11'd498, 11'd2033, 11'd344, 11'd1327, 11'd494, 11'd4270, 11'd770, 11'd4184, 11'd551, 11'd1057, 11'd3083, 11'd245, 11'd632, 11'd1222, 11'd722, 11'd107, 11'd735, 11'd1392, 11'd7, 11'd646, 11'd112, 11'd377, 11'd638, 11'd3553, 11'd78, 11'd581, 11'd65, 11'd238, 11'd2654, 11'd413, 11'd552, 11'd1954, 11'd948, 11'd500, 11'd1028, 11'd299, 11'd746, 11'd567, 11'd1328, 11'd671, 11'd310, 11'd131, 11'd89, 11'd1220, 11'd45, 11'd234, 11'd431, 11'd2110, 11'd1174, 11'd659, 11'd591, 11'd431, 11'd485, 11'd5715};

// assign sign
assign sign_o_0 = {2'd1, 2'd1, 2'd1, 2'd1, 2'd0, 2'd1, 2'd0, 2'd1, 2'd0, 2'd1, 2'd1, 2'd1, 2'd1, 2'd0, 2'd1, 2'd1, 2'd0, 2'd0, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1};
assign sign_o_1 ={2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd0, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd0, 2'd0, 2'd0, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd0, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd0, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1, 2'd1};
assign sign_o_2 = {2'd0, 2'd1, 2'd0, 2'd1, 2'd1, 2'd1, 2'd0, 2'd0, 2'd1, 2'd1, 2'd1, 2'd1, 2'd0, 2'd0, 2'd1, 2'd0, 2'd1, 2'd0, 2'd1, 2'd0, 2'd0, 2'd0, 2'd1, 2'd0, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd0, 2'd1, 2'd0, 2'd0, 2'd1, 2'd0, 2'd0, 2'd1, 2'd1, 2'd1, 2'd1, 2'd0, 2'd0, 2'd0, 2'd0, 2'd0, 2'd0, 2'd0, 2'd0, 2'd0, 2'd1, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd1, 2'd1, 2'd0, 2'd1, 2'd0, 2'd0, 2'd1, 2'd0, 2'd1};
assign sign_o_4 = {2'd1, 2'd1, 2'd0, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd1, 2'd1, 2'd1, 2'd1, 2'd0, 2'd0, 2'd0, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd1, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd1, 2'd0, 2'd0, 2'd1, 2'd1, 2'd1, 2'd1, 2'd0, 2'd1, 2'd1, 2'd1, 2'd1, 2'd0, 2'd1, 2'd0, 2'd1, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd0, 2'd0, 2'd0, 2'd0, 2'd1, 2'd1, 2'd0, 2'd1, 2'd1, 2'd0, 2'd0, 2'd1, 2'd0, 2'd1, 2'd0, 2'd0, 2'd1};

endmodule