module stimulus();

logic [0:0][27:0][27:0] test_image = {{28'b0000000000000000000000000000},{28'b0000000000000000000000000000},{28'b0000000000000000000000000000},{28'b0000000000000000000000000000},{28'b0000000000000000000000000000},{28'b0000000000000000000000000000},{28'b0000000000000000000000000000},{28'b0000000111000000000000000000},{28'b0000001111111111111110000000},{28'b0000000000111111111111000000},{28'b0000000000000000000110000000},{28'b0000000000000000000110000000},{28'b0000000000000000001100000000},{28'b0000000000000000011100000000},{28'b0000000000000000011000000000},{28'b0000000000000000111000000000},{28'b0000000000000000110000000000},{28'b0000000000000000110000000000},{28'b0000000000000001100000000000},{28'b0000000000000011100000000000},{28'b0000000000000111000000000000},{28'b0000000000000110000000000000},{28'b0000000000001100000000000000},{28'b0000000000011100000000000000},{28'b0000000000011100000000000000},{28'b0000000000011100000000000000},{28'b0000000000011000000000000000},{28'b0000000000000000000000000000}};
logic [9:0][6:0] classifier;


top bnn_test(
    .layer_i(test_image),
    .layer_o(classifier)
);

endmodule